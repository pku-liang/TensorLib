module MultiDimTime(
  input         clock,
  input         reset,
  input         io_in,
  output [1:0]  io_out_0,
  output [1:0]  io_out_1,
  output [1:0]  io_out_2,
  output [15:0] io_index_0,
  output [15:0] io_index_1,
  output [15:0] io_index_2
);
  reg [15:0] regs_0; // @[mem.scala 67:12]
  reg [31:0] _RAND_0;
  reg [15:0] regs_1; // @[mem.scala 67:12]
  reg [31:0] _RAND_1;
  reg [15:0] regs_2; // @[mem.scala 67:12]
  reg [31:0] _RAND_2;
  wire [15:0] _GEN_10 = {{15'd0}, io_in}; // @[mem.scala 69:42]
  wire [15:0] _T_1 = regs_0 + _GEN_10; // @[mem.scala 69:42]
  wire  back_0 = _T_1 == 16'hc; // @[mem.scala 69:48]
  wire [15:0] _T_3 = regs_1 + _GEN_10; // @[mem.scala 69:42]
  wire  next_1 = _T_3 == 16'h10; // @[mem.scala 69:48]
  wire [15:0] _T_5 = regs_2 + _GEN_10; // @[mem.scala 69:42]
  wire  next_2 = _T_5 == 16'h10; // @[mem.scala 69:48]
  wire  back_1 = back_0 & next_1; // @[mem.scala 71:32]
  wire  back_2 = back_1 & next_2; // @[mem.scala 71:32]
  wire  _GEN_1 = back_0 ? 1'h0 : io_in; // @[mem.scala 90:20]
  wire  _GEN_3 = back_1 ? 1'h0 : 1'h1; // @[mem.scala 79:22]
  wire  _GEN_7 = back_2 ? 1'h0 : 1'h1; // @[mem.scala 79:22]
  assign io_out_0 = {{1'd0}, _GEN_1}; // @[mem.scala 92:19 mem.scala 95:19]
  assign io_out_1 = back_0 ? {{1'd0}, _GEN_3} : 2'h2; // @[mem.scala 81:21 mem.scala 84:21 mem.scala 87:19]
  assign io_out_2 = back_1 ? {{1'd0}, _GEN_7} : 2'h2; // @[mem.scala 81:21 mem.scala 84:21 mem.scala 87:19]
  assign io_index_0 = regs_0; // @[mem.scala 76:17]
  assign io_index_1 = regs_1; // @[mem.scala 76:17]
  assign io_index_2 = regs_2; // @[mem.scala 76:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 16'h0;
    end else if (back_0) begin
      regs_0 <= 16'h0;
    end else begin
      regs_0 <= _T_1;
    end
    if (reset) begin
      regs_1 <= 16'h0;
    end else if (back_0) begin
      if (back_1) begin
        regs_1 <= 16'h0;
      end else begin
        regs_1 <= _T_3;
      end
    end
    if (reset) begin
      regs_2 <= 16'h0;
    end else if (back_1) begin
      if (back_2) begin
        regs_2 <= 16'h0;
      end else begin
        regs_2 <= _T_5;
      end
    end
  end
endmodule
module ComputeCellF(
  input          clock,
  input  [127:0] io_data_2_in_bits,
  output         io_data_2_out_valid,
  output [127:0] io_data_2_out_bits,
  input          io_data_1_in_valid,
  input  [127:0] io_data_1_in_bits,
  input          io_data_0_in_valid,
  input  [15:0]  io_data_0_in_bits
);
  wire  My_fmac_aclk; // @[cell.scala 68:62]
  wire  My_fmac_s_axis_a_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_s_axis_a_tdata; // @[cell.scala 68:62]
  wire  My_fmac_s_axis_b_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_s_axis_b_tdata; // @[cell.scala 68:62]
  wire  My_fmac_s_axis_c_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_s_axis_c_tdata; // @[cell.scala 68:62]
  wire  My_fmac_m_axis_result_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_m_axis_result_tdata; // @[cell.scala 68:62]
  wire  My_fmac_1_aclk; // @[cell.scala 68:62]
  wire  My_fmac_1_s_axis_a_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_1_s_axis_a_tdata; // @[cell.scala 68:62]
  wire  My_fmac_1_s_axis_b_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_1_s_axis_b_tdata; // @[cell.scala 68:62]
  wire  My_fmac_1_s_axis_c_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_1_s_axis_c_tdata; // @[cell.scala 68:62]
  wire  My_fmac_1_m_axis_result_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_1_m_axis_result_tdata; // @[cell.scala 68:62]
  wire  My_fmac_2_aclk; // @[cell.scala 68:62]
  wire  My_fmac_2_s_axis_a_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_2_s_axis_a_tdata; // @[cell.scala 68:62]
  wire  My_fmac_2_s_axis_b_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_2_s_axis_b_tdata; // @[cell.scala 68:62]
  wire  My_fmac_2_s_axis_c_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_2_s_axis_c_tdata; // @[cell.scala 68:62]
  wire  My_fmac_2_m_axis_result_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_2_m_axis_result_tdata; // @[cell.scala 68:62]
  wire  My_fmac_3_aclk; // @[cell.scala 68:62]
  wire  My_fmac_3_s_axis_a_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_3_s_axis_a_tdata; // @[cell.scala 68:62]
  wire  My_fmac_3_s_axis_b_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_3_s_axis_b_tdata; // @[cell.scala 68:62]
  wire  My_fmac_3_s_axis_c_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_3_s_axis_c_tdata; // @[cell.scala 68:62]
  wire  My_fmac_3_m_axis_result_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_3_m_axis_result_tdata; // @[cell.scala 68:62]
  wire  My_fmac_4_aclk; // @[cell.scala 68:62]
  wire  My_fmac_4_s_axis_a_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_4_s_axis_a_tdata; // @[cell.scala 68:62]
  wire  My_fmac_4_s_axis_b_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_4_s_axis_b_tdata; // @[cell.scala 68:62]
  wire  My_fmac_4_s_axis_c_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_4_s_axis_c_tdata; // @[cell.scala 68:62]
  wire  My_fmac_4_m_axis_result_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_4_m_axis_result_tdata; // @[cell.scala 68:62]
  wire  My_fmac_5_aclk; // @[cell.scala 68:62]
  wire  My_fmac_5_s_axis_a_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_5_s_axis_a_tdata; // @[cell.scala 68:62]
  wire  My_fmac_5_s_axis_b_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_5_s_axis_b_tdata; // @[cell.scala 68:62]
  wire  My_fmac_5_s_axis_c_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_5_s_axis_c_tdata; // @[cell.scala 68:62]
  wire  My_fmac_5_m_axis_result_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_5_m_axis_result_tdata; // @[cell.scala 68:62]
  wire  My_fmac_6_aclk; // @[cell.scala 68:62]
  wire  My_fmac_6_s_axis_a_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_6_s_axis_a_tdata; // @[cell.scala 68:62]
  wire  My_fmac_6_s_axis_b_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_6_s_axis_b_tdata; // @[cell.scala 68:62]
  wire  My_fmac_6_s_axis_c_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_6_s_axis_c_tdata; // @[cell.scala 68:62]
  wire  My_fmac_6_m_axis_result_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_6_m_axis_result_tdata; // @[cell.scala 68:62]
  wire  My_fmac_7_aclk; // @[cell.scala 68:62]
  wire  My_fmac_7_s_axis_a_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_7_s_axis_a_tdata; // @[cell.scala 68:62]
  wire  My_fmac_7_s_axis_b_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_7_s_axis_b_tdata; // @[cell.scala 68:62]
  wire  My_fmac_7_s_axis_c_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_7_s_axis_c_tdata; // @[cell.scala 68:62]
  wire  My_fmac_7_m_axis_result_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_7_m_axis_result_tdata; // @[cell.scala 68:62]
  wire [15:0] vec_b_0 = io_data_1_in_bits[15:0]; // @[cell.scala 63:35]
  wire [15:0] vec_b_1 = io_data_1_in_bits[31:16]; // @[cell.scala 63:35]
  wire [15:0] vec_b_2 = io_data_1_in_bits[47:32]; // @[cell.scala 63:35]
  wire [15:0] vec_b_3 = io_data_1_in_bits[63:48]; // @[cell.scala 63:35]
  wire [15:0] vec_b_4 = io_data_1_in_bits[79:64]; // @[cell.scala 63:35]
  wire [15:0] vec_b_5 = io_data_1_in_bits[95:80]; // @[cell.scala 63:35]
  wire [15:0] vec_b_6 = io_data_1_in_bits[111:96]; // @[cell.scala 63:35]
  wire [15:0] vec_b_7 = io_data_1_in_bits[127:112]; // @[cell.scala 63:35]
  wire [15:0] vec_c_in_0 = io_data_2_in_bits[15:0]; // @[cell.scala 66:38]
  wire [15:0] vec_c_in_1 = io_data_2_in_bits[31:16]; // @[cell.scala 66:38]
  wire [15:0] vec_c_in_2 = io_data_2_in_bits[47:32]; // @[cell.scala 66:38]
  wire [15:0] vec_c_in_3 = io_data_2_in_bits[63:48]; // @[cell.scala 66:38]
  wire [15:0] vec_c_in_4 = io_data_2_in_bits[79:64]; // @[cell.scala 66:38]
  wire [15:0] vec_c_in_5 = io_data_2_in_bits[95:80]; // @[cell.scala 66:38]
  wire [15:0] vec_c_in_6 = io_data_2_in_bits[111:96]; // @[cell.scala 66:38]
  wire [15:0] vec_c_in_7 = io_data_2_in_bits[127:112]; // @[cell.scala 66:38]
  wire [15:0] vec_c_out_1 = My_fmac_1_m_axis_result_tdata[15:0]; // @[cell.scala 58:25 cell.scala 88:30]
  wire [15:0] vec_c_out_0 = My_fmac_m_axis_result_tdata[15:0]; // @[cell.scala 58:25 cell.scala 88:30]
  wire [15:0] vec_c_out_3 = My_fmac_3_m_axis_result_tdata[15:0]; // @[cell.scala 58:25 cell.scala 88:30]
  wire [15:0] vec_c_out_2 = My_fmac_2_m_axis_result_tdata[15:0]; // @[cell.scala 58:25 cell.scala 88:30]
  wire [63:0] _T_22 = {vec_c_out_3,vec_c_out_2,vec_c_out_1,vec_c_out_0}; // @[cell.scala 91:38]
  wire [15:0] vec_c_out_5 = My_fmac_5_m_axis_result_tdata[15:0]; // @[cell.scala 58:25 cell.scala 88:30]
  wire [15:0] vec_c_out_4 = My_fmac_4_m_axis_result_tdata[15:0]; // @[cell.scala 58:25 cell.scala 88:30]
  wire [15:0] vec_c_out_7 = My_fmac_7_m_axis_result_tdata[15:0]; // @[cell.scala 58:25 cell.scala 88:30]
  wire [15:0] vec_c_out_6 = My_fmac_6_m_axis_result_tdata[15:0]; // @[cell.scala 58:25 cell.scala 88:30]
  wire [63:0] _T_25 = {vec_c_out_7,vec_c_out_6,vec_c_out_5,vec_c_out_4}; // @[cell.scala 91:38]
  My_fmac My_fmac ( // @[cell.scala 68:62]
    .aclk(My_fmac_aclk),
    .s_axis_a_tvalid(My_fmac_s_axis_a_tvalid),
    .s_axis_a_tdata(My_fmac_s_axis_a_tdata),
    .s_axis_b_tvalid(My_fmac_s_axis_b_tvalid),
    .s_axis_b_tdata(My_fmac_s_axis_b_tdata),
    .s_axis_c_tvalid(My_fmac_s_axis_c_tvalid),
    .s_axis_c_tdata(My_fmac_s_axis_c_tdata),
    .m_axis_result_tvalid(My_fmac_m_axis_result_tvalid),
    .m_axis_result_tdata(My_fmac_m_axis_result_tdata)
  );
  My_fmac My_fmac_1 ( // @[cell.scala 68:62]
    .aclk(My_fmac_1_aclk),
    .s_axis_a_tvalid(My_fmac_1_s_axis_a_tvalid),
    .s_axis_a_tdata(My_fmac_1_s_axis_a_tdata),
    .s_axis_b_tvalid(My_fmac_1_s_axis_b_tvalid),
    .s_axis_b_tdata(My_fmac_1_s_axis_b_tdata),
    .s_axis_c_tvalid(My_fmac_1_s_axis_c_tvalid),
    .s_axis_c_tdata(My_fmac_1_s_axis_c_tdata),
    .m_axis_result_tvalid(My_fmac_1_m_axis_result_tvalid),
    .m_axis_result_tdata(My_fmac_1_m_axis_result_tdata)
  );
  My_fmac My_fmac_2 ( // @[cell.scala 68:62]
    .aclk(My_fmac_2_aclk),
    .s_axis_a_tvalid(My_fmac_2_s_axis_a_tvalid),
    .s_axis_a_tdata(My_fmac_2_s_axis_a_tdata),
    .s_axis_b_tvalid(My_fmac_2_s_axis_b_tvalid),
    .s_axis_b_tdata(My_fmac_2_s_axis_b_tdata),
    .s_axis_c_tvalid(My_fmac_2_s_axis_c_tvalid),
    .s_axis_c_tdata(My_fmac_2_s_axis_c_tdata),
    .m_axis_result_tvalid(My_fmac_2_m_axis_result_tvalid),
    .m_axis_result_tdata(My_fmac_2_m_axis_result_tdata)
  );
  My_fmac My_fmac_3 ( // @[cell.scala 68:62]
    .aclk(My_fmac_3_aclk),
    .s_axis_a_tvalid(My_fmac_3_s_axis_a_tvalid),
    .s_axis_a_tdata(My_fmac_3_s_axis_a_tdata),
    .s_axis_b_tvalid(My_fmac_3_s_axis_b_tvalid),
    .s_axis_b_tdata(My_fmac_3_s_axis_b_tdata),
    .s_axis_c_tvalid(My_fmac_3_s_axis_c_tvalid),
    .s_axis_c_tdata(My_fmac_3_s_axis_c_tdata),
    .m_axis_result_tvalid(My_fmac_3_m_axis_result_tvalid),
    .m_axis_result_tdata(My_fmac_3_m_axis_result_tdata)
  );
  My_fmac My_fmac_4 ( // @[cell.scala 68:62]
    .aclk(My_fmac_4_aclk),
    .s_axis_a_tvalid(My_fmac_4_s_axis_a_tvalid),
    .s_axis_a_tdata(My_fmac_4_s_axis_a_tdata),
    .s_axis_b_tvalid(My_fmac_4_s_axis_b_tvalid),
    .s_axis_b_tdata(My_fmac_4_s_axis_b_tdata),
    .s_axis_c_tvalid(My_fmac_4_s_axis_c_tvalid),
    .s_axis_c_tdata(My_fmac_4_s_axis_c_tdata),
    .m_axis_result_tvalid(My_fmac_4_m_axis_result_tvalid),
    .m_axis_result_tdata(My_fmac_4_m_axis_result_tdata)
  );
  My_fmac My_fmac_5 ( // @[cell.scala 68:62]
    .aclk(My_fmac_5_aclk),
    .s_axis_a_tvalid(My_fmac_5_s_axis_a_tvalid),
    .s_axis_a_tdata(My_fmac_5_s_axis_a_tdata),
    .s_axis_b_tvalid(My_fmac_5_s_axis_b_tvalid),
    .s_axis_b_tdata(My_fmac_5_s_axis_b_tdata),
    .s_axis_c_tvalid(My_fmac_5_s_axis_c_tvalid),
    .s_axis_c_tdata(My_fmac_5_s_axis_c_tdata),
    .m_axis_result_tvalid(My_fmac_5_m_axis_result_tvalid),
    .m_axis_result_tdata(My_fmac_5_m_axis_result_tdata)
  );
  My_fmac My_fmac_6 ( // @[cell.scala 68:62]
    .aclk(My_fmac_6_aclk),
    .s_axis_a_tvalid(My_fmac_6_s_axis_a_tvalid),
    .s_axis_a_tdata(My_fmac_6_s_axis_a_tdata),
    .s_axis_b_tvalid(My_fmac_6_s_axis_b_tvalid),
    .s_axis_b_tdata(My_fmac_6_s_axis_b_tdata),
    .s_axis_c_tvalid(My_fmac_6_s_axis_c_tvalid),
    .s_axis_c_tdata(My_fmac_6_s_axis_c_tdata),
    .m_axis_result_tvalid(My_fmac_6_m_axis_result_tvalid),
    .m_axis_result_tdata(My_fmac_6_m_axis_result_tdata)
  );
  My_fmac My_fmac_7 ( // @[cell.scala 68:62]
    .aclk(My_fmac_7_aclk),
    .s_axis_a_tvalid(My_fmac_7_s_axis_a_tvalid),
    .s_axis_a_tdata(My_fmac_7_s_axis_a_tdata),
    .s_axis_b_tvalid(My_fmac_7_s_axis_b_tvalid),
    .s_axis_b_tdata(My_fmac_7_s_axis_b_tdata),
    .s_axis_c_tvalid(My_fmac_7_s_axis_c_tvalid),
    .s_axis_c_tdata(My_fmac_7_s_axis_c_tdata),
    .m_axis_result_tvalid(My_fmac_7_m_axis_result_tvalid),
    .m_axis_result_tdata(My_fmac_7_m_axis_result_tdata)
  );
  assign io_data_2_out_valid = My_fmac_m_axis_result_tvalid; // @[cell.scala 94:26]
  assign io_data_2_out_bits = {_T_25,_T_22}; // @[cell.scala 91:25]
  assign My_fmac_aclk = clock; // @[cell.scala 81:31]
  assign My_fmac_s_axis_a_tvalid = io_data_0_in_valid; // @[cell.scala 82:41]
  assign My_fmac_s_axis_a_tdata = {{16'd0}, io_data_0_in_bits}; // @[cell.scala 84:40]
  assign My_fmac_s_axis_b_tvalid = io_data_1_in_valid; // @[cell.scala 83:41]
  assign My_fmac_s_axis_b_tdata = {{16'd0}, vec_b_0}; // @[cell.scala 85:40]
  assign My_fmac_s_axis_c_tvalid = 1'h1; // @[cell.scala 86:41]
  assign My_fmac_s_axis_c_tdata = {{16'd0}, vec_c_in_0}; // @[cell.scala 87:40]
  assign My_fmac_1_aclk = clock; // @[cell.scala 81:31]
  assign My_fmac_1_s_axis_a_tvalid = io_data_0_in_valid; // @[cell.scala 82:41]
  assign My_fmac_1_s_axis_a_tdata = {{16'd0}, io_data_0_in_bits}; // @[cell.scala 84:40]
  assign My_fmac_1_s_axis_b_tvalid = io_data_1_in_valid; // @[cell.scala 83:41]
  assign My_fmac_1_s_axis_b_tdata = {{16'd0}, vec_b_1}; // @[cell.scala 85:40]
  assign My_fmac_1_s_axis_c_tvalid = 1'h1; // @[cell.scala 86:41]
  assign My_fmac_1_s_axis_c_tdata = {{16'd0}, vec_c_in_1}; // @[cell.scala 87:40]
  assign My_fmac_2_aclk = clock; // @[cell.scala 81:31]
  assign My_fmac_2_s_axis_a_tvalid = io_data_0_in_valid; // @[cell.scala 82:41]
  assign My_fmac_2_s_axis_a_tdata = {{16'd0}, io_data_0_in_bits}; // @[cell.scala 84:40]
  assign My_fmac_2_s_axis_b_tvalid = io_data_1_in_valid; // @[cell.scala 83:41]
  assign My_fmac_2_s_axis_b_tdata = {{16'd0}, vec_b_2}; // @[cell.scala 85:40]
  assign My_fmac_2_s_axis_c_tvalid = 1'h1; // @[cell.scala 86:41]
  assign My_fmac_2_s_axis_c_tdata = {{16'd0}, vec_c_in_2}; // @[cell.scala 87:40]
  assign My_fmac_3_aclk = clock; // @[cell.scala 81:31]
  assign My_fmac_3_s_axis_a_tvalid = io_data_0_in_valid; // @[cell.scala 82:41]
  assign My_fmac_3_s_axis_a_tdata = {{16'd0}, io_data_0_in_bits}; // @[cell.scala 84:40]
  assign My_fmac_3_s_axis_b_tvalid = io_data_1_in_valid; // @[cell.scala 83:41]
  assign My_fmac_3_s_axis_b_tdata = {{16'd0}, vec_b_3}; // @[cell.scala 85:40]
  assign My_fmac_3_s_axis_c_tvalid = 1'h1; // @[cell.scala 86:41]
  assign My_fmac_3_s_axis_c_tdata = {{16'd0}, vec_c_in_3}; // @[cell.scala 87:40]
  assign My_fmac_4_aclk = clock; // @[cell.scala 81:31]
  assign My_fmac_4_s_axis_a_tvalid = io_data_0_in_valid; // @[cell.scala 82:41]
  assign My_fmac_4_s_axis_a_tdata = {{16'd0}, io_data_0_in_bits}; // @[cell.scala 84:40]
  assign My_fmac_4_s_axis_b_tvalid = io_data_1_in_valid; // @[cell.scala 83:41]
  assign My_fmac_4_s_axis_b_tdata = {{16'd0}, vec_b_4}; // @[cell.scala 85:40]
  assign My_fmac_4_s_axis_c_tvalid = 1'h1; // @[cell.scala 86:41]
  assign My_fmac_4_s_axis_c_tdata = {{16'd0}, vec_c_in_4}; // @[cell.scala 87:40]
  assign My_fmac_5_aclk = clock; // @[cell.scala 81:31]
  assign My_fmac_5_s_axis_a_tvalid = io_data_0_in_valid; // @[cell.scala 82:41]
  assign My_fmac_5_s_axis_a_tdata = {{16'd0}, io_data_0_in_bits}; // @[cell.scala 84:40]
  assign My_fmac_5_s_axis_b_tvalid = io_data_1_in_valid; // @[cell.scala 83:41]
  assign My_fmac_5_s_axis_b_tdata = {{16'd0}, vec_b_5}; // @[cell.scala 85:40]
  assign My_fmac_5_s_axis_c_tvalid = 1'h1; // @[cell.scala 86:41]
  assign My_fmac_5_s_axis_c_tdata = {{16'd0}, vec_c_in_5}; // @[cell.scala 87:40]
  assign My_fmac_6_aclk = clock; // @[cell.scala 81:31]
  assign My_fmac_6_s_axis_a_tvalid = io_data_0_in_valid; // @[cell.scala 82:41]
  assign My_fmac_6_s_axis_a_tdata = {{16'd0}, io_data_0_in_bits}; // @[cell.scala 84:40]
  assign My_fmac_6_s_axis_b_tvalid = io_data_1_in_valid; // @[cell.scala 83:41]
  assign My_fmac_6_s_axis_b_tdata = {{16'd0}, vec_b_6}; // @[cell.scala 85:40]
  assign My_fmac_6_s_axis_c_tvalid = 1'h1; // @[cell.scala 86:41]
  assign My_fmac_6_s_axis_c_tdata = {{16'd0}, vec_c_in_6}; // @[cell.scala 87:40]
  assign My_fmac_7_aclk = clock; // @[cell.scala 81:31]
  assign My_fmac_7_s_axis_a_tvalid = io_data_0_in_valid; // @[cell.scala 82:41]
  assign My_fmac_7_s_axis_a_tdata = {{16'd0}, io_data_0_in_bits}; // @[cell.scala 84:40]
  assign My_fmac_7_s_axis_b_tvalid = io_data_1_in_valid; // @[cell.scala 83:41]
  assign My_fmac_7_s_axis_b_tdata = {{16'd0}, vec_b_7}; // @[cell.scala 85:40]
  assign My_fmac_7_s_axis_c_tvalid = 1'h1; // @[cell.scala 86:41]
  assign My_fmac_7_s_axis_c_tdata = {{16'd0}, vec_c_in_7}; // @[cell.scala 87:40]
endmodule
module SystolicInput(
  input         clock,
  input         reset,
  input         io_port_in_valid,
  input  [15:0] io_port_in_bits,
  output        io_port_out_valid,
  output [15:0] io_port_out_bits,
  output        io_to_cell_valid,
  output [15:0] io_to_cell_bits
);
  reg [15:0] reg_bits; // @[pe_modules.scala 55:18]
  reg [31:0] _RAND_0;
  reg  reg_valid; // @[pe_modules.scala 55:18]
  reg [31:0] _RAND_1;
  reg [15:0] to_cell_delay1_bits; // @[pe_modules.scala 55:18]
  reg [31:0] _RAND_2;
  reg  to_cell_delay1_valid; // @[pe_modules.scala 55:18]
  reg [31:0] _RAND_3;
  reg [15:0] to_cell_delay2_bits; // @[pe_modules.scala 55:18]
  reg [31:0] _RAND_4;
  reg  to_cell_delay2_valid; // @[pe_modules.scala 55:18]
  reg [31:0] _RAND_5;
  assign io_port_out_valid = reg_valid; // @[pe_modules.scala 87:15]
  assign io_port_out_bits = reg_bits; // @[pe_modules.scala 87:15]
  assign io_to_cell_valid = to_cell_delay2_valid; // @[pe_modules.scala 88:14]
  assign io_to_cell_bits = to_cell_delay2_bits; // @[pe_modules.scala 88:14]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_bits = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  reg_valid = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  to_cell_delay1_bits = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  to_cell_delay1_valid = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  to_cell_delay2_bits = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  to_cell_delay2_valid = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      reg_bits <= 16'h0;
    end else begin
      reg_bits <= io_port_in_bits;
    end
    if (reset) begin
      reg_valid <= 1'h0;
    end else begin
      reg_valid <= io_port_in_valid;
    end
    if (reset) begin
      to_cell_delay1_bits <= 16'h0;
    end else begin
      to_cell_delay1_bits <= reg_bits;
    end
    if (reset) begin
      to_cell_delay1_valid <= 1'h0;
    end else begin
      to_cell_delay1_valid <= reg_valid;
    end
    if (reset) begin
      to_cell_delay2_bits <= 16'h0;
    end else begin
      to_cell_delay2_bits <= to_cell_delay1_bits;
    end
    if (reset) begin
      to_cell_delay2_valid <= 1'h0;
    end else begin
      to_cell_delay2_valid <= to_cell_delay1_valid;
    end
  end
endmodule
module SystolicInput_1(
  input          clock,
  input          reset,
  input          io_port_in_valid,
  input  [127:0] io_port_in_bits,
  output         io_port_out_valid,
  output [127:0] io_port_out_bits,
  output         io_to_cell_valid,
  output [127:0] io_to_cell_bits
);
  reg [127:0] reg_bits; // @[pe_modules.scala 55:18]
  reg [127:0] _RAND_0;
  reg  reg_valid; // @[pe_modules.scala 55:18]
  reg [31:0] _RAND_1;
  reg [127:0] to_cell_delay1_bits; // @[pe_modules.scala 55:18]
  reg [127:0] _RAND_2;
  reg  to_cell_delay1_valid; // @[pe_modules.scala 55:18]
  reg [31:0] _RAND_3;
  reg [127:0] to_cell_delay2_bits; // @[pe_modules.scala 55:18]
  reg [127:0] _RAND_4;
  reg  to_cell_delay2_valid; // @[pe_modules.scala 55:18]
  reg [31:0] _RAND_5;
  assign io_port_out_valid = reg_valid; // @[pe_modules.scala 87:15]
  assign io_port_out_bits = reg_bits; // @[pe_modules.scala 87:15]
  assign io_to_cell_valid = to_cell_delay2_valid; // @[pe_modules.scala 88:14]
  assign io_to_cell_bits = to_cell_delay2_bits; // @[pe_modules.scala 88:14]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {4{`RANDOM}};
  reg_bits = _RAND_0[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  reg_valid = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {4{`RANDOM}};
  to_cell_delay1_bits = _RAND_2[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  to_cell_delay1_valid = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {4{`RANDOM}};
  to_cell_delay2_bits = _RAND_4[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  to_cell_delay2_valid = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      reg_bits <= 128'h0;
    end else begin
      reg_bits <= io_port_in_bits;
    end
    if (reset) begin
      reg_valid <= 1'h0;
    end else begin
      reg_valid <= io_port_in_valid;
    end
    if (reset) begin
      to_cell_delay1_bits <= 128'h0;
    end else begin
      to_cell_delay1_bits <= reg_bits;
    end
    if (reset) begin
      to_cell_delay1_valid <= 1'h0;
    end else begin
      to_cell_delay1_valid <= reg_valid;
    end
    if (reset) begin
      to_cell_delay2_bits <= 128'h0;
    end else begin
      to_cell_delay2_bits <= to_cell_delay1_bits;
    end
    if (reset) begin
      to_cell_delay2_valid <= 1'h0;
    end else begin
      to_cell_delay2_valid <= to_cell_delay1_valid;
    end
  end
endmodule
module StationaryOutput_OutCell(
  input          clock,
  input          reset,
  output         io_port_out_valid,
  output [127:0] io_port_out_bits,
  input          io_port_sig_stat2trans,
  input          io_from_cell_valid,
  input  [127:0] io_from_cell_bits,
  output [127:0] io_to_cell_bits
);
  reg  reg_stat2trans; // @[pe_modules.scala 161:31]
  reg [31:0] _RAND_0;
  assign io_port_out_valid = reg_stat2trans & io_from_cell_valid; // @[pe_modules.scala 167:23 pe_modules.scala 171:23]
  assign io_port_out_bits = reg_stat2trans ? io_from_cell_bits : 128'h0; // @[pe_modules.scala 166:22 pe_modules.scala 170:22]
  assign io_to_cell_bits = reg_stat2trans ? 128'h0 : io_from_cell_bits; // @[pe_modules.scala 174:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_stat2trans = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      reg_stat2trans <= 1'h0;
    end else begin
      reg_stat2trans <= io_port_sig_stat2trans;
    end
  end
endmodule
module PE(
  input          clock,
  input          reset,
  output         io_data_2_out_valid,
  output [127:0] io_data_2_out_bits,
  input          io_data_2_sig_stat2trans,
  input          io_data_1_in_valid,
  input  [127:0] io_data_1_in_bits,
  output         io_data_1_out_valid,
  output [127:0] io_data_1_out_bits,
  input          io_data_0_in_valid,
  input  [15:0]  io_data_0_in_bits,
  output         io_data_0_out_valid,
  output [15:0]  io_data_0_out_bits
);
  wire  ComputeCellF_clock; // @[pe.scala 44:11]
  wire [127:0] ComputeCellF_io_data_2_in_bits; // @[pe.scala 44:11]
  wire  ComputeCellF_io_data_2_out_valid; // @[pe.scala 44:11]
  wire [127:0] ComputeCellF_io_data_2_out_bits; // @[pe.scala 44:11]
  wire  ComputeCellF_io_data_1_in_valid; // @[pe.scala 44:11]
  wire [127:0] ComputeCellF_io_data_1_in_bits; // @[pe.scala 44:11]
  wire  ComputeCellF_io_data_0_in_valid; // @[pe.scala 44:11]
  wire [15:0] ComputeCellF_io_data_0_in_bits; // @[pe.scala 44:11]
  wire  SystolicInput_clock; // @[pe.scala 46:11]
  wire  SystolicInput_reset; // @[pe.scala 46:11]
  wire  SystolicInput_io_port_in_valid; // @[pe.scala 46:11]
  wire [15:0] SystolicInput_io_port_in_bits; // @[pe.scala 46:11]
  wire  SystolicInput_io_port_out_valid; // @[pe.scala 46:11]
  wire [15:0] SystolicInput_io_port_out_bits; // @[pe.scala 46:11]
  wire  SystolicInput_io_to_cell_valid; // @[pe.scala 46:11]
  wire [15:0] SystolicInput_io_to_cell_bits; // @[pe.scala 46:11]
  wire  SystolicInput_1_clock; // @[pe.scala 46:11]
  wire  SystolicInput_1_reset; // @[pe.scala 46:11]
  wire  SystolicInput_1_io_port_in_valid; // @[pe.scala 46:11]
  wire [127:0] SystolicInput_1_io_port_in_bits; // @[pe.scala 46:11]
  wire  SystolicInput_1_io_port_out_valid; // @[pe.scala 46:11]
  wire [127:0] SystolicInput_1_io_port_out_bits; // @[pe.scala 46:11]
  wire  SystolicInput_1_io_to_cell_valid; // @[pe.scala 46:11]
  wire [127:0] SystolicInput_1_io_to_cell_bits; // @[pe.scala 46:11]
  wire  StationaryOutput_OutCell_clock; // @[pe.scala 46:11]
  wire  StationaryOutput_OutCell_reset; // @[pe.scala 46:11]
  wire  StationaryOutput_OutCell_io_port_out_valid; // @[pe.scala 46:11]
  wire [127:0] StationaryOutput_OutCell_io_port_out_bits; // @[pe.scala 46:11]
  wire  StationaryOutput_OutCell_io_port_sig_stat2trans; // @[pe.scala 46:11]
  wire  StationaryOutput_OutCell_io_from_cell_valid; // @[pe.scala 46:11]
  wire [127:0] StationaryOutput_OutCell_io_from_cell_bits; // @[pe.scala 46:11]
  wire [127:0] StationaryOutput_OutCell_io_to_cell_bits; // @[pe.scala 46:11]
  ComputeCellF ComputeCellF ( // @[pe.scala 44:11]
    .clock(ComputeCellF_clock),
    .io_data_2_in_bits(ComputeCellF_io_data_2_in_bits),
    .io_data_2_out_valid(ComputeCellF_io_data_2_out_valid),
    .io_data_2_out_bits(ComputeCellF_io_data_2_out_bits),
    .io_data_1_in_valid(ComputeCellF_io_data_1_in_valid),
    .io_data_1_in_bits(ComputeCellF_io_data_1_in_bits),
    .io_data_0_in_valid(ComputeCellF_io_data_0_in_valid),
    .io_data_0_in_bits(ComputeCellF_io_data_0_in_bits)
  );
  SystolicInput SystolicInput ( // @[pe.scala 46:11]
    .clock(SystolicInput_clock),
    .reset(SystolicInput_reset),
    .io_port_in_valid(SystolicInput_io_port_in_valid),
    .io_port_in_bits(SystolicInput_io_port_in_bits),
    .io_port_out_valid(SystolicInput_io_port_out_valid),
    .io_port_out_bits(SystolicInput_io_port_out_bits),
    .io_to_cell_valid(SystolicInput_io_to_cell_valid),
    .io_to_cell_bits(SystolicInput_io_to_cell_bits)
  );
  SystolicInput_1 SystolicInput_1 ( // @[pe.scala 46:11]
    .clock(SystolicInput_1_clock),
    .reset(SystolicInput_1_reset),
    .io_port_in_valid(SystolicInput_1_io_port_in_valid),
    .io_port_in_bits(SystolicInput_1_io_port_in_bits),
    .io_port_out_valid(SystolicInput_1_io_port_out_valid),
    .io_port_out_bits(SystolicInput_1_io_port_out_bits),
    .io_to_cell_valid(SystolicInput_1_io_to_cell_valid),
    .io_to_cell_bits(SystolicInput_1_io_to_cell_bits)
  );
  StationaryOutput_OutCell StationaryOutput_OutCell ( // @[pe.scala 46:11]
    .clock(StationaryOutput_OutCell_clock),
    .reset(StationaryOutput_OutCell_reset),
    .io_port_out_valid(StationaryOutput_OutCell_io_port_out_valid),
    .io_port_out_bits(StationaryOutput_OutCell_io_port_out_bits),
    .io_port_sig_stat2trans(StationaryOutput_OutCell_io_port_sig_stat2trans),
    .io_from_cell_valid(StationaryOutput_OutCell_io_from_cell_valid),
    .io_from_cell_bits(StationaryOutput_OutCell_io_from_cell_bits),
    .io_to_cell_bits(StationaryOutput_OutCell_io_to_cell_bits)
  );
  assign io_data_2_out_valid = StationaryOutput_OutCell_io_port_out_valid; // @[pe.scala 52:20]
  assign io_data_2_out_bits = StationaryOutput_OutCell_io_port_out_bits; // @[pe.scala 52:20]
  assign io_data_1_out_valid = SystolicInput_1_io_port_out_valid; // @[pe.scala 52:20]
  assign io_data_1_out_bits = SystolicInput_1_io_port_out_bits; // @[pe.scala 52:20]
  assign io_data_0_out_valid = SystolicInput_io_port_out_valid; // @[pe.scala 52:20]
  assign io_data_0_out_bits = SystolicInput_io_port_out_bits; // @[pe.scala 52:20]
  assign ComputeCellF_clock = clock;
  assign ComputeCellF_io_data_2_in_bits = StationaryOutput_OutCell_io_to_cell_bits; // @[pe.scala 53:19]
  assign ComputeCellF_io_data_1_in_valid = SystolicInput_1_io_to_cell_valid; // @[pe.scala 53:19]
  assign ComputeCellF_io_data_1_in_bits = SystolicInput_1_io_to_cell_bits; // @[pe.scala 53:19]
  assign ComputeCellF_io_data_0_in_valid = SystolicInput_io_to_cell_valid; // @[pe.scala 53:19]
  assign ComputeCellF_io_data_0_in_bits = SystolicInput_io_to_cell_bits; // @[pe.scala 53:19]
  assign SystolicInput_clock = clock;
  assign SystolicInput_reset = reset;
  assign SystolicInput_io_port_in_valid = io_data_0_in_valid; // @[pe.scala 51:20]
  assign SystolicInput_io_port_in_bits = io_data_0_in_bits; // @[pe.scala 51:20]
  assign SystolicInput_1_clock = clock;
  assign SystolicInput_1_reset = reset;
  assign SystolicInput_1_io_port_in_valid = io_data_1_in_valid; // @[pe.scala 51:20]
  assign SystolicInput_1_io_port_in_bits = io_data_1_in_bits; // @[pe.scala 51:20]
  assign StationaryOutput_OutCell_clock = clock;
  assign StationaryOutput_OutCell_reset = reset;
  assign StationaryOutput_OutCell_io_port_sig_stat2trans = io_data_2_sig_stat2trans; // @[pe.scala 64:38]
  assign StationaryOutput_OutCell_io_from_cell_valid = ComputeCellF_io_data_2_out_valid; // @[pe.scala 57:28]
  assign StationaryOutput_OutCell_io_from_cell_bits = ComputeCellF_io_data_2_out_bits; // @[pe.scala 57:28]
endmodule
module PENetwork(
  output        io_to_pes_0_in_valid,
  output [15:0] io_to_pes_0_in_bits,
  input         io_to_pes_0_out_valid,
  input  [15:0] io_to_pes_0_out_bits,
  output        io_to_pes_1_in_valid,
  output [15:0] io_to_pes_1_in_bits,
  input         io_to_pes_1_out_valid,
  input  [15:0] io_to_pes_1_out_bits,
  output        io_to_pes_2_in_valid,
  output [15:0] io_to_pes_2_in_bits,
  input         io_to_pes_2_out_valid,
  input  [15:0] io_to_pes_2_out_bits,
  output        io_to_pes_3_in_valid,
  output [15:0] io_to_pes_3_in_bits,
  input         io_to_pes_3_out_valid,
  input  [15:0] io_to_pes_3_out_bits,
  output        io_to_pes_4_in_valid,
  output [15:0] io_to_pes_4_in_bits,
  input         io_to_pes_4_out_valid,
  input  [15:0] io_to_pes_4_out_bits,
  output        io_to_pes_5_in_valid,
  output [15:0] io_to_pes_5_in_bits,
  input         io_to_pes_5_out_valid,
  input  [15:0] io_to_pes_5_out_bits,
  output        io_to_pes_6_in_valid,
  output [15:0] io_to_pes_6_in_bits,
  input         io_to_pes_6_out_valid,
  input  [15:0] io_to_pes_6_out_bits,
  output        io_to_pes_7_in_valid,
  output [15:0] io_to_pes_7_in_bits,
  input         io_to_pes_7_out_valid,
  input  [15:0] io_to_pes_7_out_bits,
  output        io_to_pes_8_in_valid,
  output [15:0] io_to_pes_8_in_bits,
  input         io_to_pes_8_out_valid,
  input  [15:0] io_to_pes_8_out_bits,
  output        io_to_pes_9_in_valid,
  output [15:0] io_to_pes_9_in_bits,
  input         io_to_pes_9_out_valid,
  input  [15:0] io_to_pes_9_out_bits,
  output        io_to_pes_10_in_valid,
  output [15:0] io_to_pes_10_in_bits,
  input         io_to_pes_10_out_valid,
  input  [15:0] io_to_pes_10_out_bits,
  output        io_to_pes_11_in_valid,
  output [15:0] io_to_pes_11_in_bits,
  input         io_to_pes_11_out_valid,
  input  [15:0] io_to_pes_11_out_bits,
  output        io_to_pes_12_in_valid,
  output [15:0] io_to_pes_12_in_bits,
  input         io_to_pes_12_out_valid,
  input  [15:0] io_to_pes_12_out_bits,
  output        io_to_pes_13_in_valid,
  output [15:0] io_to_pes_13_in_bits,
  input         io_to_pes_13_out_valid,
  input  [15:0] io_to_pes_13_out_bits,
  output        io_to_pes_14_in_valid,
  output [15:0] io_to_pes_14_in_bits,
  input         io_to_pes_14_out_valid,
  input  [15:0] io_to_pes_14_out_bits,
  output        io_to_pes_15_in_valid,
  output [15:0] io_to_pes_15_in_bits,
  input         io_to_pes_15_out_valid,
  input  [15:0] io_to_pes_15_out_bits,
  output        io_to_pes_16_in_valid,
  output [15:0] io_to_pes_16_in_bits,
  input         io_to_pes_16_out_valid,
  input  [15:0] io_to_pes_16_out_bits,
  output        io_to_pes_17_in_valid,
  output [15:0] io_to_pes_17_in_bits,
  input         io_to_pes_17_out_valid,
  input  [15:0] io_to_pes_17_out_bits,
  output        io_to_pes_18_in_valid,
  output [15:0] io_to_pes_18_in_bits,
  input         io_to_pes_18_out_valid,
  input  [15:0] io_to_pes_18_out_bits,
  output        io_to_pes_19_in_valid,
  output [15:0] io_to_pes_19_in_bits,
  input         io_to_pes_19_out_valid,
  input  [15:0] io_to_pes_19_out_bits,
  output        io_to_pes_20_in_valid,
  output [15:0] io_to_pes_20_in_bits,
  input         io_to_pes_20_out_valid,
  input  [15:0] io_to_pes_20_out_bits,
  output        io_to_pes_21_in_valid,
  output [15:0] io_to_pes_21_in_bits,
  input         io_to_pes_21_out_valid,
  input  [15:0] io_to_pes_21_out_bits,
  output        io_to_pes_22_in_valid,
  output [15:0] io_to_pes_22_in_bits,
  input         io_to_pes_22_out_valid,
  input  [15:0] io_to_pes_22_out_bits,
  output        io_to_pes_23_in_valid,
  output [15:0] io_to_pes_23_in_bits,
  input         io_to_pes_23_out_valid,
  input  [15:0] io_to_pes_23_out_bits,
  output        io_to_pes_24_in_valid,
  output [15:0] io_to_pes_24_in_bits,
  input         io_to_pes_24_out_valid,
  input  [15:0] io_to_pes_24_out_bits,
  output        io_to_pes_25_in_valid,
  output [15:0] io_to_pes_25_in_bits,
  input         io_to_pes_25_out_valid,
  input  [15:0] io_to_pes_25_out_bits,
  output        io_to_pes_26_in_valid,
  output [15:0] io_to_pes_26_in_bits,
  input         io_to_pes_26_out_valid,
  input  [15:0] io_to_pes_26_out_bits,
  output        io_to_pes_27_in_valid,
  output [15:0] io_to_pes_27_in_bits,
  input         io_to_pes_27_out_valid,
  input  [15:0] io_to_pes_27_out_bits,
  output        io_to_pes_28_in_valid,
  output [15:0] io_to_pes_28_in_bits,
  input         io_to_pes_28_out_valid,
  input  [15:0] io_to_pes_28_out_bits,
  output        io_to_pes_29_in_valid,
  output [15:0] io_to_pes_29_in_bits,
  input         io_to_mem_valid,
  input  [15:0] io_to_mem_bits
);
  assign io_to_pes_0_in_valid = io_to_mem_valid; // @[pe.scala 128:23]
  assign io_to_pes_0_in_bits = io_to_mem_bits; // @[pe.scala 128:23]
  assign io_to_pes_1_in_valid = io_to_pes_0_out_valid; // @[pe.scala 125:23]
  assign io_to_pes_1_in_bits = io_to_pes_0_out_bits; // @[pe.scala 125:23]
  assign io_to_pes_2_in_valid = io_to_pes_1_out_valid; // @[pe.scala 125:23]
  assign io_to_pes_2_in_bits = io_to_pes_1_out_bits; // @[pe.scala 125:23]
  assign io_to_pes_3_in_valid = io_to_pes_2_out_valid; // @[pe.scala 125:23]
  assign io_to_pes_3_in_bits = io_to_pes_2_out_bits; // @[pe.scala 125:23]
  assign io_to_pes_4_in_valid = io_to_pes_3_out_valid; // @[pe.scala 125:23]
  assign io_to_pes_4_in_bits = io_to_pes_3_out_bits; // @[pe.scala 125:23]
  assign io_to_pes_5_in_valid = io_to_pes_4_out_valid; // @[pe.scala 125:23]
  assign io_to_pes_5_in_bits = io_to_pes_4_out_bits; // @[pe.scala 125:23]
  assign io_to_pes_6_in_valid = io_to_pes_5_out_valid; // @[pe.scala 125:23]
  assign io_to_pes_6_in_bits = io_to_pes_5_out_bits; // @[pe.scala 125:23]
  assign io_to_pes_7_in_valid = io_to_pes_6_out_valid; // @[pe.scala 125:23]
  assign io_to_pes_7_in_bits = io_to_pes_6_out_bits; // @[pe.scala 125:23]
  assign io_to_pes_8_in_valid = io_to_pes_7_out_valid; // @[pe.scala 125:23]
  assign io_to_pes_8_in_bits = io_to_pes_7_out_bits; // @[pe.scala 125:23]
  assign io_to_pes_9_in_valid = io_to_pes_8_out_valid; // @[pe.scala 125:23]
  assign io_to_pes_9_in_bits = io_to_pes_8_out_bits; // @[pe.scala 125:23]
  assign io_to_pes_10_in_valid = io_to_pes_9_out_valid; // @[pe.scala 125:23]
  assign io_to_pes_10_in_bits = io_to_pes_9_out_bits; // @[pe.scala 125:23]
  assign io_to_pes_11_in_valid = io_to_pes_10_out_valid; // @[pe.scala 125:23]
  assign io_to_pes_11_in_bits = io_to_pes_10_out_bits; // @[pe.scala 125:23]
  assign io_to_pes_12_in_valid = io_to_pes_11_out_valid; // @[pe.scala 125:23]
  assign io_to_pes_12_in_bits = io_to_pes_11_out_bits; // @[pe.scala 125:23]
  assign io_to_pes_13_in_valid = io_to_pes_12_out_valid; // @[pe.scala 125:23]
  assign io_to_pes_13_in_bits = io_to_pes_12_out_bits; // @[pe.scala 125:23]
  assign io_to_pes_14_in_valid = io_to_pes_13_out_valid; // @[pe.scala 125:23]
  assign io_to_pes_14_in_bits = io_to_pes_13_out_bits; // @[pe.scala 125:23]
  assign io_to_pes_15_in_valid = io_to_pes_14_out_valid; // @[pe.scala 125:23]
  assign io_to_pes_15_in_bits = io_to_pes_14_out_bits; // @[pe.scala 125:23]
  assign io_to_pes_16_in_valid = io_to_pes_15_out_valid; // @[pe.scala 125:23]
  assign io_to_pes_16_in_bits = io_to_pes_15_out_bits; // @[pe.scala 125:23]
  assign io_to_pes_17_in_valid = io_to_pes_16_out_valid; // @[pe.scala 125:23]
  assign io_to_pes_17_in_bits = io_to_pes_16_out_bits; // @[pe.scala 125:23]
  assign io_to_pes_18_in_valid = io_to_pes_17_out_valid; // @[pe.scala 125:23]
  assign io_to_pes_18_in_bits = io_to_pes_17_out_bits; // @[pe.scala 125:23]
  assign io_to_pes_19_in_valid = io_to_pes_18_out_valid; // @[pe.scala 125:23]
  assign io_to_pes_19_in_bits = io_to_pes_18_out_bits; // @[pe.scala 125:23]
  assign io_to_pes_20_in_valid = io_to_pes_19_out_valid; // @[pe.scala 125:23]
  assign io_to_pes_20_in_bits = io_to_pes_19_out_bits; // @[pe.scala 125:23]
  assign io_to_pes_21_in_valid = io_to_pes_20_out_valid; // @[pe.scala 125:23]
  assign io_to_pes_21_in_bits = io_to_pes_20_out_bits; // @[pe.scala 125:23]
  assign io_to_pes_22_in_valid = io_to_pes_21_out_valid; // @[pe.scala 125:23]
  assign io_to_pes_22_in_bits = io_to_pes_21_out_bits; // @[pe.scala 125:23]
  assign io_to_pes_23_in_valid = io_to_pes_22_out_valid; // @[pe.scala 125:23]
  assign io_to_pes_23_in_bits = io_to_pes_22_out_bits; // @[pe.scala 125:23]
  assign io_to_pes_24_in_valid = io_to_pes_23_out_valid; // @[pe.scala 125:23]
  assign io_to_pes_24_in_bits = io_to_pes_23_out_bits; // @[pe.scala 125:23]
  assign io_to_pes_25_in_valid = io_to_pes_24_out_valid; // @[pe.scala 125:23]
  assign io_to_pes_25_in_bits = io_to_pes_24_out_bits; // @[pe.scala 125:23]
  assign io_to_pes_26_in_valid = io_to_pes_25_out_valid; // @[pe.scala 125:23]
  assign io_to_pes_26_in_bits = io_to_pes_25_out_bits; // @[pe.scala 125:23]
  assign io_to_pes_27_in_valid = io_to_pes_26_out_valid; // @[pe.scala 125:23]
  assign io_to_pes_27_in_bits = io_to_pes_26_out_bits; // @[pe.scala 125:23]
  assign io_to_pes_28_in_valid = io_to_pes_27_out_valid; // @[pe.scala 125:23]
  assign io_to_pes_28_in_bits = io_to_pes_27_out_bits; // @[pe.scala 125:23]
  assign io_to_pes_29_in_valid = io_to_pes_28_out_valid; // @[pe.scala 125:23]
  assign io_to_pes_29_in_bits = io_to_pes_28_out_bits; // @[pe.scala 125:23]
endmodule
module PENetwork_22(
  output         io_to_pes_0_in_valid,
  output [127:0] io_to_pes_0_in_bits,
  input          io_to_pes_0_out_valid,
  input  [127:0] io_to_pes_0_out_bits,
  output         io_to_pes_1_in_valid,
  output [127:0] io_to_pes_1_in_bits,
  input          io_to_pes_1_out_valid,
  input  [127:0] io_to_pes_1_out_bits,
  output         io_to_pes_2_in_valid,
  output [127:0] io_to_pes_2_in_bits,
  input          io_to_pes_2_out_valid,
  input  [127:0] io_to_pes_2_out_bits,
  output         io_to_pes_3_in_valid,
  output [127:0] io_to_pes_3_in_bits,
  input          io_to_pes_3_out_valid,
  input  [127:0] io_to_pes_3_out_bits,
  output         io_to_pes_4_in_valid,
  output [127:0] io_to_pes_4_in_bits,
  input          io_to_pes_4_out_valid,
  input  [127:0] io_to_pes_4_out_bits,
  output         io_to_pes_5_in_valid,
  output [127:0] io_to_pes_5_in_bits,
  input          io_to_pes_5_out_valid,
  input  [127:0] io_to_pes_5_out_bits,
  output         io_to_pes_6_in_valid,
  output [127:0] io_to_pes_6_in_bits,
  input          io_to_pes_6_out_valid,
  input  [127:0] io_to_pes_6_out_bits,
  output         io_to_pes_7_in_valid,
  output [127:0] io_to_pes_7_in_bits,
  input          io_to_pes_7_out_valid,
  input  [127:0] io_to_pes_7_out_bits,
  output         io_to_pes_8_in_valid,
  output [127:0] io_to_pes_8_in_bits,
  input          io_to_pes_8_out_valid,
  input  [127:0] io_to_pes_8_out_bits,
  output         io_to_pes_9_in_valid,
  output [127:0] io_to_pes_9_in_bits,
  input          io_to_pes_9_out_valid,
  input  [127:0] io_to_pes_9_out_bits,
  output         io_to_pes_10_in_valid,
  output [127:0] io_to_pes_10_in_bits,
  input          io_to_pes_10_out_valid,
  input  [127:0] io_to_pes_10_out_bits,
  output         io_to_pes_11_in_valid,
  output [127:0] io_to_pes_11_in_bits,
  input          io_to_pes_11_out_valid,
  input  [127:0] io_to_pes_11_out_bits,
  output         io_to_pes_12_in_valid,
  output [127:0] io_to_pes_12_in_bits,
  input          io_to_pes_12_out_valid,
  input  [127:0] io_to_pes_12_out_bits,
  output         io_to_pes_13_in_valid,
  output [127:0] io_to_pes_13_in_bits,
  input          io_to_pes_13_out_valid,
  input  [127:0] io_to_pes_13_out_bits,
  output         io_to_pes_14_in_valid,
  output [127:0] io_to_pes_14_in_bits,
  input          io_to_pes_14_out_valid,
  input  [127:0] io_to_pes_14_out_bits,
  output         io_to_pes_15_in_valid,
  output [127:0] io_to_pes_15_in_bits,
  input          io_to_pes_15_out_valid,
  input  [127:0] io_to_pes_15_out_bits,
  output         io_to_pes_16_in_valid,
  output [127:0] io_to_pes_16_in_bits,
  input          io_to_pes_16_out_valid,
  input  [127:0] io_to_pes_16_out_bits,
  output         io_to_pes_17_in_valid,
  output [127:0] io_to_pes_17_in_bits,
  input          io_to_pes_17_out_valid,
  input  [127:0] io_to_pes_17_out_bits,
  output         io_to_pes_18_in_valid,
  output [127:0] io_to_pes_18_in_bits,
  input          io_to_pes_18_out_valid,
  input  [127:0] io_to_pes_18_out_bits,
  output         io_to_pes_19_in_valid,
  output [127:0] io_to_pes_19_in_bits,
  input          io_to_pes_19_out_valid,
  input  [127:0] io_to_pes_19_out_bits,
  output         io_to_pes_20_in_valid,
  output [127:0] io_to_pes_20_in_bits,
  input          io_to_pes_20_out_valid,
  input  [127:0] io_to_pes_20_out_bits,
  output         io_to_pes_21_in_valid,
  output [127:0] io_to_pes_21_in_bits,
  input          io_to_mem_valid,
  input  [127:0] io_to_mem_bits
);
  assign io_to_pes_0_in_valid = io_to_mem_valid; // @[pe.scala 128:23]
  assign io_to_pes_0_in_bits = io_to_mem_bits; // @[pe.scala 128:23]
  assign io_to_pes_1_in_valid = io_to_pes_0_out_valid; // @[pe.scala 125:23]
  assign io_to_pes_1_in_bits = io_to_pes_0_out_bits; // @[pe.scala 125:23]
  assign io_to_pes_2_in_valid = io_to_pes_1_out_valid; // @[pe.scala 125:23]
  assign io_to_pes_2_in_bits = io_to_pes_1_out_bits; // @[pe.scala 125:23]
  assign io_to_pes_3_in_valid = io_to_pes_2_out_valid; // @[pe.scala 125:23]
  assign io_to_pes_3_in_bits = io_to_pes_2_out_bits; // @[pe.scala 125:23]
  assign io_to_pes_4_in_valid = io_to_pes_3_out_valid; // @[pe.scala 125:23]
  assign io_to_pes_4_in_bits = io_to_pes_3_out_bits; // @[pe.scala 125:23]
  assign io_to_pes_5_in_valid = io_to_pes_4_out_valid; // @[pe.scala 125:23]
  assign io_to_pes_5_in_bits = io_to_pes_4_out_bits; // @[pe.scala 125:23]
  assign io_to_pes_6_in_valid = io_to_pes_5_out_valid; // @[pe.scala 125:23]
  assign io_to_pes_6_in_bits = io_to_pes_5_out_bits; // @[pe.scala 125:23]
  assign io_to_pes_7_in_valid = io_to_pes_6_out_valid; // @[pe.scala 125:23]
  assign io_to_pes_7_in_bits = io_to_pes_6_out_bits; // @[pe.scala 125:23]
  assign io_to_pes_8_in_valid = io_to_pes_7_out_valid; // @[pe.scala 125:23]
  assign io_to_pes_8_in_bits = io_to_pes_7_out_bits; // @[pe.scala 125:23]
  assign io_to_pes_9_in_valid = io_to_pes_8_out_valid; // @[pe.scala 125:23]
  assign io_to_pes_9_in_bits = io_to_pes_8_out_bits; // @[pe.scala 125:23]
  assign io_to_pes_10_in_valid = io_to_pes_9_out_valid; // @[pe.scala 125:23]
  assign io_to_pes_10_in_bits = io_to_pes_9_out_bits; // @[pe.scala 125:23]
  assign io_to_pes_11_in_valid = io_to_pes_10_out_valid; // @[pe.scala 125:23]
  assign io_to_pes_11_in_bits = io_to_pes_10_out_bits; // @[pe.scala 125:23]
  assign io_to_pes_12_in_valid = io_to_pes_11_out_valid; // @[pe.scala 125:23]
  assign io_to_pes_12_in_bits = io_to_pes_11_out_bits; // @[pe.scala 125:23]
  assign io_to_pes_13_in_valid = io_to_pes_12_out_valid; // @[pe.scala 125:23]
  assign io_to_pes_13_in_bits = io_to_pes_12_out_bits; // @[pe.scala 125:23]
  assign io_to_pes_14_in_valid = io_to_pes_13_out_valid; // @[pe.scala 125:23]
  assign io_to_pes_14_in_bits = io_to_pes_13_out_bits; // @[pe.scala 125:23]
  assign io_to_pes_15_in_valid = io_to_pes_14_out_valid; // @[pe.scala 125:23]
  assign io_to_pes_15_in_bits = io_to_pes_14_out_bits; // @[pe.scala 125:23]
  assign io_to_pes_16_in_valid = io_to_pes_15_out_valid; // @[pe.scala 125:23]
  assign io_to_pes_16_in_bits = io_to_pes_15_out_bits; // @[pe.scala 125:23]
  assign io_to_pes_17_in_valid = io_to_pes_16_out_valid; // @[pe.scala 125:23]
  assign io_to_pes_17_in_bits = io_to_pes_16_out_bits; // @[pe.scala 125:23]
  assign io_to_pes_18_in_valid = io_to_pes_17_out_valid; // @[pe.scala 125:23]
  assign io_to_pes_18_in_bits = io_to_pes_17_out_bits; // @[pe.scala 125:23]
  assign io_to_pes_19_in_valid = io_to_pes_18_out_valid; // @[pe.scala 125:23]
  assign io_to_pes_19_in_bits = io_to_pes_18_out_bits; // @[pe.scala 125:23]
  assign io_to_pes_20_in_valid = io_to_pes_19_out_valid; // @[pe.scala 125:23]
  assign io_to_pes_20_in_bits = io_to_pes_19_out_bits; // @[pe.scala 125:23]
  assign io_to_pes_21_in_valid = io_to_pes_20_out_valid; // @[pe.scala 125:23]
  assign io_to_pes_21_in_bits = io_to_pes_20_out_bits; // @[pe.scala 125:23]
endmodule
module PENetwork_52(
  input          clock,
  input          reset,
  input          io_to_pes_0_out_valid,
  input  [127:0] io_to_pes_0_out_bits,
  output         io_to_pes_0_sig_stat2trans,
  input          io_to_pes_1_out_valid,
  input  [127:0] io_to_pes_1_out_bits,
  output         io_to_pes_1_sig_stat2trans,
  input          io_to_pes_2_out_valid,
  input  [127:0] io_to_pes_2_out_bits,
  output         io_to_pes_2_sig_stat2trans,
  input          io_to_pes_3_out_valid,
  input  [127:0] io_to_pes_3_out_bits,
  output         io_to_pes_3_sig_stat2trans,
  input          io_to_pes_4_out_valid,
  input  [127:0] io_to_pes_4_out_bits,
  output         io_to_pes_4_sig_stat2trans,
  input          io_to_pes_5_out_valid,
  input  [127:0] io_to_pes_5_out_bits,
  output         io_to_pes_5_sig_stat2trans,
  input          io_to_pes_6_out_valid,
  input  [127:0] io_to_pes_6_out_bits,
  output         io_to_pes_6_sig_stat2trans,
  input          io_to_pes_7_out_valid,
  input  [127:0] io_to_pes_7_out_bits,
  output         io_to_pes_7_sig_stat2trans,
  input          io_to_pes_8_out_valid,
  input  [127:0] io_to_pes_8_out_bits,
  output         io_to_pes_8_sig_stat2trans,
  input          io_to_pes_9_out_valid,
  input  [127:0] io_to_pes_9_out_bits,
  output         io_to_pes_9_sig_stat2trans,
  input          io_to_pes_10_out_valid,
  input  [127:0] io_to_pes_10_out_bits,
  output         io_to_pes_10_sig_stat2trans,
  input          io_to_pes_11_out_valid,
  input  [127:0] io_to_pes_11_out_bits,
  output         io_to_pes_11_sig_stat2trans,
  input          io_to_pes_12_out_valid,
  input  [127:0] io_to_pes_12_out_bits,
  output         io_to_pes_12_sig_stat2trans,
  input          io_to_pes_13_out_valid,
  input  [127:0] io_to_pes_13_out_bits,
  output         io_to_pes_13_sig_stat2trans,
  input          io_to_pes_14_out_valid,
  input  [127:0] io_to_pes_14_out_bits,
  output         io_to_pes_14_sig_stat2trans,
  input          io_to_pes_15_out_valid,
  input  [127:0] io_to_pes_15_out_bits,
  output         io_to_pes_15_sig_stat2trans,
  input          io_to_pes_16_out_valid,
  input  [127:0] io_to_pes_16_out_bits,
  output         io_to_pes_16_sig_stat2trans,
  input          io_to_pes_17_out_valid,
  input  [127:0] io_to_pes_17_out_bits,
  output         io_to_pes_17_sig_stat2trans,
  input          io_to_pes_18_out_valid,
  input  [127:0] io_to_pes_18_out_bits,
  output         io_to_pes_18_sig_stat2trans,
  input          io_to_pes_19_out_valid,
  input  [127:0] io_to_pes_19_out_bits,
  output         io_to_pes_19_sig_stat2trans,
  input          io_to_pes_20_out_valid,
  input  [127:0] io_to_pes_20_out_bits,
  output         io_to_pes_20_sig_stat2trans,
  input          io_to_pes_21_out_valid,
  input  [127:0] io_to_pes_21_out_bits,
  output         io_to_pes_21_sig_stat2trans,
  output         io_to_mem_valid,
  output [127:0] io_to_mem_bits,
  input          io_sig_stat2trans
);
  reg [127:0] _T [0:11]; // @[pe.scala 94:49]
  reg [127:0] _RAND_0;
  wire [127:0] _T__T_195_data; // @[pe.scala 94:49]
  wire [3:0] _T__T_195_addr; // @[pe.scala 94:49]
  reg [127:0] _RAND_1;
  wire [127:0] _T__T_48_data; // @[pe.scala 94:49]
  wire [3:0] _T__T_48_addr; // @[pe.scala 94:49]
  wire  _T__T_48_mask; // @[pe.scala 94:49]
  wire  _T__T_48_en; // @[pe.scala 94:49]
  reg  _T__T_195_en_pipe_0;
  reg [31:0] _RAND_2;
  reg [3:0] _T__T_195_addr_pipe_0;
  reg [31:0] _RAND_3;
  reg [127:0] _T_1 [0:11]; // @[pe.scala 94:49]
  reg [127:0] _RAND_4;
  wire [127:0] _T_1__T_197_data; // @[pe.scala 94:49]
  wire [3:0] _T_1__T_197_addr; // @[pe.scala 94:49]
  reg [127:0] _RAND_5;
  wire [127:0] _T_1__T_54_data; // @[pe.scala 94:49]
  wire [3:0] _T_1__T_54_addr; // @[pe.scala 94:49]
  wire  _T_1__T_54_mask; // @[pe.scala 94:49]
  wire  _T_1__T_54_en; // @[pe.scala 94:49]
  reg  _T_1__T_197_en_pipe_0;
  reg [31:0] _RAND_6;
  reg [3:0] _T_1__T_197_addr_pipe_0;
  reg [31:0] _RAND_7;
  reg [127:0] _T_2 [0:11]; // @[pe.scala 94:49]
  reg [127:0] _RAND_8;
  wire [127:0] _T_2__T_199_data; // @[pe.scala 94:49]
  wire [3:0] _T_2__T_199_addr; // @[pe.scala 94:49]
  reg [127:0] _RAND_9;
  wire [127:0] _T_2__T_60_data; // @[pe.scala 94:49]
  wire [3:0] _T_2__T_60_addr; // @[pe.scala 94:49]
  wire  _T_2__T_60_mask; // @[pe.scala 94:49]
  wire  _T_2__T_60_en; // @[pe.scala 94:49]
  reg  _T_2__T_199_en_pipe_0;
  reg [31:0] _RAND_10;
  reg [3:0] _T_2__T_199_addr_pipe_0;
  reg [31:0] _RAND_11;
  reg [127:0] _T_3 [0:11]; // @[pe.scala 94:49]
  reg [127:0] _RAND_12;
  wire [127:0] _T_3__T_201_data; // @[pe.scala 94:49]
  wire [3:0] _T_3__T_201_addr; // @[pe.scala 94:49]
  reg [127:0] _RAND_13;
  wire [127:0] _T_3__T_66_data; // @[pe.scala 94:49]
  wire [3:0] _T_3__T_66_addr; // @[pe.scala 94:49]
  wire  _T_3__T_66_mask; // @[pe.scala 94:49]
  wire  _T_3__T_66_en; // @[pe.scala 94:49]
  reg  _T_3__T_201_en_pipe_0;
  reg [31:0] _RAND_14;
  reg [3:0] _T_3__T_201_addr_pipe_0;
  reg [31:0] _RAND_15;
  reg [127:0] _T_4 [0:11]; // @[pe.scala 94:49]
  reg [127:0] _RAND_16;
  wire [127:0] _T_4__T_203_data; // @[pe.scala 94:49]
  wire [3:0] _T_4__T_203_addr; // @[pe.scala 94:49]
  reg [127:0] _RAND_17;
  wire [127:0] _T_4__T_72_data; // @[pe.scala 94:49]
  wire [3:0] _T_4__T_72_addr; // @[pe.scala 94:49]
  wire  _T_4__T_72_mask; // @[pe.scala 94:49]
  wire  _T_4__T_72_en; // @[pe.scala 94:49]
  reg  _T_4__T_203_en_pipe_0;
  reg [31:0] _RAND_18;
  reg [3:0] _T_4__T_203_addr_pipe_0;
  reg [31:0] _RAND_19;
  reg [127:0] _T_5 [0:11]; // @[pe.scala 94:49]
  reg [127:0] _RAND_20;
  wire [127:0] _T_5__T_205_data; // @[pe.scala 94:49]
  wire [3:0] _T_5__T_205_addr; // @[pe.scala 94:49]
  reg [127:0] _RAND_21;
  wire [127:0] _T_5__T_78_data; // @[pe.scala 94:49]
  wire [3:0] _T_5__T_78_addr; // @[pe.scala 94:49]
  wire  _T_5__T_78_mask; // @[pe.scala 94:49]
  wire  _T_5__T_78_en; // @[pe.scala 94:49]
  reg  _T_5__T_205_en_pipe_0;
  reg [31:0] _RAND_22;
  reg [3:0] _T_5__T_205_addr_pipe_0;
  reg [31:0] _RAND_23;
  reg [127:0] _T_6 [0:11]; // @[pe.scala 94:49]
  reg [127:0] _RAND_24;
  wire [127:0] _T_6__T_207_data; // @[pe.scala 94:49]
  wire [3:0] _T_6__T_207_addr; // @[pe.scala 94:49]
  reg [127:0] _RAND_25;
  wire [127:0] _T_6__T_84_data; // @[pe.scala 94:49]
  wire [3:0] _T_6__T_84_addr; // @[pe.scala 94:49]
  wire  _T_6__T_84_mask; // @[pe.scala 94:49]
  wire  _T_6__T_84_en; // @[pe.scala 94:49]
  reg  _T_6__T_207_en_pipe_0;
  reg [31:0] _RAND_26;
  reg [3:0] _T_6__T_207_addr_pipe_0;
  reg [31:0] _RAND_27;
  reg [127:0] _T_7 [0:11]; // @[pe.scala 94:49]
  reg [127:0] _RAND_28;
  wire [127:0] _T_7__T_209_data; // @[pe.scala 94:49]
  wire [3:0] _T_7__T_209_addr; // @[pe.scala 94:49]
  reg [127:0] _RAND_29;
  wire [127:0] _T_7__T_90_data; // @[pe.scala 94:49]
  wire [3:0] _T_7__T_90_addr; // @[pe.scala 94:49]
  wire  _T_7__T_90_mask; // @[pe.scala 94:49]
  wire  _T_7__T_90_en; // @[pe.scala 94:49]
  reg  _T_7__T_209_en_pipe_0;
  reg [31:0] _RAND_30;
  reg [3:0] _T_7__T_209_addr_pipe_0;
  reg [31:0] _RAND_31;
  reg [127:0] _T_8 [0:11]; // @[pe.scala 94:49]
  reg [127:0] _RAND_32;
  wire [127:0] _T_8__T_211_data; // @[pe.scala 94:49]
  wire [3:0] _T_8__T_211_addr; // @[pe.scala 94:49]
  reg [127:0] _RAND_33;
  wire [127:0] _T_8__T_96_data; // @[pe.scala 94:49]
  wire [3:0] _T_8__T_96_addr; // @[pe.scala 94:49]
  wire  _T_8__T_96_mask; // @[pe.scala 94:49]
  wire  _T_8__T_96_en; // @[pe.scala 94:49]
  reg  _T_8__T_211_en_pipe_0;
  reg [31:0] _RAND_34;
  reg [3:0] _T_8__T_211_addr_pipe_0;
  reg [31:0] _RAND_35;
  reg [127:0] _T_9 [0:11]; // @[pe.scala 94:49]
  reg [127:0] _RAND_36;
  wire [127:0] _T_9__T_213_data; // @[pe.scala 94:49]
  wire [3:0] _T_9__T_213_addr; // @[pe.scala 94:49]
  reg [127:0] _RAND_37;
  wire [127:0] _T_9__T_102_data; // @[pe.scala 94:49]
  wire [3:0] _T_9__T_102_addr; // @[pe.scala 94:49]
  wire  _T_9__T_102_mask; // @[pe.scala 94:49]
  wire  _T_9__T_102_en; // @[pe.scala 94:49]
  reg  _T_9__T_213_en_pipe_0;
  reg [31:0] _RAND_38;
  reg [3:0] _T_9__T_213_addr_pipe_0;
  reg [31:0] _RAND_39;
  reg [127:0] _T_10 [0:11]; // @[pe.scala 94:49]
  reg [127:0] _RAND_40;
  wire [127:0] _T_10__T_215_data; // @[pe.scala 94:49]
  wire [3:0] _T_10__T_215_addr; // @[pe.scala 94:49]
  reg [127:0] _RAND_41;
  wire [127:0] _T_10__T_108_data; // @[pe.scala 94:49]
  wire [3:0] _T_10__T_108_addr; // @[pe.scala 94:49]
  wire  _T_10__T_108_mask; // @[pe.scala 94:49]
  wire  _T_10__T_108_en; // @[pe.scala 94:49]
  reg  _T_10__T_215_en_pipe_0;
  reg [31:0] _RAND_42;
  reg [3:0] _T_10__T_215_addr_pipe_0;
  reg [31:0] _RAND_43;
  reg [127:0] _T_11 [0:11]; // @[pe.scala 94:49]
  reg [127:0] _RAND_44;
  wire [127:0] _T_11__T_217_data; // @[pe.scala 94:49]
  wire [3:0] _T_11__T_217_addr; // @[pe.scala 94:49]
  reg [127:0] _RAND_45;
  wire [127:0] _T_11__T_114_data; // @[pe.scala 94:49]
  wire [3:0] _T_11__T_114_addr; // @[pe.scala 94:49]
  wire  _T_11__T_114_mask; // @[pe.scala 94:49]
  wire  _T_11__T_114_en; // @[pe.scala 94:49]
  reg  _T_11__T_217_en_pipe_0;
  reg [31:0] _RAND_46;
  reg [3:0] _T_11__T_217_addr_pipe_0;
  reg [31:0] _RAND_47;
  reg [127:0] _T_12 [0:11]; // @[pe.scala 94:49]
  reg [127:0] _RAND_48;
  wire [127:0] _T_12__T_219_data; // @[pe.scala 94:49]
  wire [3:0] _T_12__T_219_addr; // @[pe.scala 94:49]
  reg [127:0] _RAND_49;
  wire [127:0] _T_12__T_120_data; // @[pe.scala 94:49]
  wire [3:0] _T_12__T_120_addr; // @[pe.scala 94:49]
  wire  _T_12__T_120_mask; // @[pe.scala 94:49]
  wire  _T_12__T_120_en; // @[pe.scala 94:49]
  reg  _T_12__T_219_en_pipe_0;
  reg [31:0] _RAND_50;
  reg [3:0] _T_12__T_219_addr_pipe_0;
  reg [31:0] _RAND_51;
  reg [127:0] _T_13 [0:11]; // @[pe.scala 94:49]
  reg [127:0] _RAND_52;
  wire [127:0] _T_13__T_221_data; // @[pe.scala 94:49]
  wire [3:0] _T_13__T_221_addr; // @[pe.scala 94:49]
  reg [127:0] _RAND_53;
  wire [127:0] _T_13__T_126_data; // @[pe.scala 94:49]
  wire [3:0] _T_13__T_126_addr; // @[pe.scala 94:49]
  wire  _T_13__T_126_mask; // @[pe.scala 94:49]
  wire  _T_13__T_126_en; // @[pe.scala 94:49]
  reg  _T_13__T_221_en_pipe_0;
  reg [31:0] _RAND_54;
  reg [3:0] _T_13__T_221_addr_pipe_0;
  reg [31:0] _RAND_55;
  reg [127:0] _T_14 [0:11]; // @[pe.scala 94:49]
  reg [127:0] _RAND_56;
  wire [127:0] _T_14__T_223_data; // @[pe.scala 94:49]
  wire [3:0] _T_14__T_223_addr; // @[pe.scala 94:49]
  reg [127:0] _RAND_57;
  wire [127:0] _T_14__T_132_data; // @[pe.scala 94:49]
  wire [3:0] _T_14__T_132_addr; // @[pe.scala 94:49]
  wire  _T_14__T_132_mask; // @[pe.scala 94:49]
  wire  _T_14__T_132_en; // @[pe.scala 94:49]
  reg  _T_14__T_223_en_pipe_0;
  reg [31:0] _RAND_58;
  reg [3:0] _T_14__T_223_addr_pipe_0;
  reg [31:0] _RAND_59;
  reg [127:0] _T_15 [0:11]; // @[pe.scala 94:49]
  reg [127:0] _RAND_60;
  wire [127:0] _T_15__T_225_data; // @[pe.scala 94:49]
  wire [3:0] _T_15__T_225_addr; // @[pe.scala 94:49]
  reg [127:0] _RAND_61;
  wire [127:0] _T_15__T_138_data; // @[pe.scala 94:49]
  wire [3:0] _T_15__T_138_addr; // @[pe.scala 94:49]
  wire  _T_15__T_138_mask; // @[pe.scala 94:49]
  wire  _T_15__T_138_en; // @[pe.scala 94:49]
  reg  _T_15__T_225_en_pipe_0;
  reg [31:0] _RAND_62;
  reg [3:0] _T_15__T_225_addr_pipe_0;
  reg [31:0] _RAND_63;
  reg [127:0] _T_16 [0:11]; // @[pe.scala 94:49]
  reg [127:0] _RAND_64;
  wire [127:0] _T_16__T_227_data; // @[pe.scala 94:49]
  wire [3:0] _T_16__T_227_addr; // @[pe.scala 94:49]
  reg [127:0] _RAND_65;
  wire [127:0] _T_16__T_144_data; // @[pe.scala 94:49]
  wire [3:0] _T_16__T_144_addr; // @[pe.scala 94:49]
  wire  _T_16__T_144_mask; // @[pe.scala 94:49]
  wire  _T_16__T_144_en; // @[pe.scala 94:49]
  reg  _T_16__T_227_en_pipe_0;
  reg [31:0] _RAND_66;
  reg [3:0] _T_16__T_227_addr_pipe_0;
  reg [31:0] _RAND_67;
  reg [127:0] _T_17 [0:11]; // @[pe.scala 94:49]
  reg [127:0] _RAND_68;
  wire [127:0] _T_17__T_229_data; // @[pe.scala 94:49]
  wire [3:0] _T_17__T_229_addr; // @[pe.scala 94:49]
  reg [127:0] _RAND_69;
  wire [127:0] _T_17__T_150_data; // @[pe.scala 94:49]
  wire [3:0] _T_17__T_150_addr; // @[pe.scala 94:49]
  wire  _T_17__T_150_mask; // @[pe.scala 94:49]
  wire  _T_17__T_150_en; // @[pe.scala 94:49]
  reg  _T_17__T_229_en_pipe_0;
  reg [31:0] _RAND_70;
  reg [3:0] _T_17__T_229_addr_pipe_0;
  reg [31:0] _RAND_71;
  reg [127:0] _T_18 [0:11]; // @[pe.scala 94:49]
  reg [127:0] _RAND_72;
  wire [127:0] _T_18__T_231_data; // @[pe.scala 94:49]
  wire [3:0] _T_18__T_231_addr; // @[pe.scala 94:49]
  reg [127:0] _RAND_73;
  wire [127:0] _T_18__T_156_data; // @[pe.scala 94:49]
  wire [3:0] _T_18__T_156_addr; // @[pe.scala 94:49]
  wire  _T_18__T_156_mask; // @[pe.scala 94:49]
  wire  _T_18__T_156_en; // @[pe.scala 94:49]
  reg  _T_18__T_231_en_pipe_0;
  reg [31:0] _RAND_74;
  reg [3:0] _T_18__T_231_addr_pipe_0;
  reg [31:0] _RAND_75;
  reg [127:0] _T_19 [0:11]; // @[pe.scala 94:49]
  reg [127:0] _RAND_76;
  wire [127:0] _T_19__T_233_data; // @[pe.scala 94:49]
  wire [3:0] _T_19__T_233_addr; // @[pe.scala 94:49]
  reg [127:0] _RAND_77;
  wire [127:0] _T_19__T_162_data; // @[pe.scala 94:49]
  wire [3:0] _T_19__T_162_addr; // @[pe.scala 94:49]
  wire  _T_19__T_162_mask; // @[pe.scala 94:49]
  wire  _T_19__T_162_en; // @[pe.scala 94:49]
  reg  _T_19__T_233_en_pipe_0;
  reg [31:0] _RAND_78;
  reg [3:0] _T_19__T_233_addr_pipe_0;
  reg [31:0] _RAND_79;
  reg [127:0] _T_20 [0:11]; // @[pe.scala 94:49]
  reg [127:0] _RAND_80;
  wire [127:0] _T_20__T_235_data; // @[pe.scala 94:49]
  wire [3:0] _T_20__T_235_addr; // @[pe.scala 94:49]
  reg [127:0] _RAND_81;
  wire [127:0] _T_20__T_168_data; // @[pe.scala 94:49]
  wire [3:0] _T_20__T_168_addr; // @[pe.scala 94:49]
  wire  _T_20__T_168_mask; // @[pe.scala 94:49]
  wire  _T_20__T_168_en; // @[pe.scala 94:49]
  reg  _T_20__T_235_en_pipe_0;
  reg [31:0] _RAND_82;
  reg [3:0] _T_20__T_235_addr_pipe_0;
  reg [31:0] _RAND_83;
  reg [127:0] _T_21 [0:11]; // @[pe.scala 94:49]
  reg [127:0] _RAND_84;
  wire [127:0] _T_21__T_237_data; // @[pe.scala 94:49]
  wire [3:0] _T_21__T_237_addr; // @[pe.scala 94:49]
  reg [127:0] _RAND_85;
  wire [127:0] _T_21__T_174_data; // @[pe.scala 94:49]
  wire [3:0] _T_21__T_174_addr; // @[pe.scala 94:49]
  wire  _T_21__T_174_mask; // @[pe.scala 94:49]
  wire  _T_21__T_174_en; // @[pe.scala 94:49]
  reg  _T_21__T_237_en_pipe_0;
  reg [31:0] _RAND_86;
  reg [3:0] _T_21__T_237_addr_pipe_0;
  reg [31:0] _RAND_87;
  reg [4:0] _T_22; // @[pe.scala 95:44]
  reg [31:0] _RAND_88;
  reg [4:0] _T_23; // @[pe.scala 95:44]
  reg [31:0] _RAND_89;
  reg [4:0] _T_24; // @[pe.scala 95:44]
  reg [31:0] _RAND_90;
  reg [4:0] _T_25; // @[pe.scala 95:44]
  reg [31:0] _RAND_91;
  reg [4:0] _T_26; // @[pe.scala 95:44]
  reg [31:0] _RAND_92;
  reg [4:0] _T_27; // @[pe.scala 95:44]
  reg [31:0] _RAND_93;
  reg [4:0] _T_28; // @[pe.scala 95:44]
  reg [31:0] _RAND_94;
  reg [4:0] _T_29; // @[pe.scala 95:44]
  reg [31:0] _RAND_95;
  reg [4:0] _T_30; // @[pe.scala 95:44]
  reg [31:0] _RAND_96;
  reg [4:0] _T_31; // @[pe.scala 95:44]
  reg [31:0] _RAND_97;
  reg [4:0] _T_32; // @[pe.scala 95:44]
  reg [31:0] _RAND_98;
  reg [4:0] _T_33; // @[pe.scala 95:44]
  reg [31:0] _RAND_99;
  reg [4:0] _T_34; // @[pe.scala 95:44]
  reg [31:0] _RAND_100;
  reg [4:0] _T_35; // @[pe.scala 95:44]
  reg [31:0] _RAND_101;
  reg [4:0] _T_36; // @[pe.scala 95:44]
  reg [31:0] _RAND_102;
  reg [4:0] _T_37; // @[pe.scala 95:44]
  reg [31:0] _RAND_103;
  reg [4:0] _T_38; // @[pe.scala 95:44]
  reg [31:0] _RAND_104;
  reg [4:0] _T_39; // @[pe.scala 95:44]
  reg [31:0] _RAND_105;
  reg [4:0] _T_40; // @[pe.scala 95:44]
  reg [31:0] _RAND_106;
  reg [4:0] _T_41; // @[pe.scala 95:44]
  reg [31:0] _RAND_107;
  reg [4:0] _T_42; // @[pe.scala 95:44]
  reg [31:0] _RAND_108;
  reg [4:0] _T_43; // @[pe.scala 95:44]
  reg [31:0] _RAND_109;
  reg  _T_44; // @[pe.scala 96:29]
  reg [31:0] _RAND_110;
  reg [9:0] _T_45; // @[pe.scala 97:26]
  reg [31:0] _RAND_111;
  reg [9:0] _T_46; // @[pe.scala 98:25]
  reg [31:0] _RAND_112;
  wire  _T_49 = _T_22 == 5'hb; // @[pe.scala 106:35]
  wire [4:0] _T_51 = _T_22 + 5'h1; // @[pe.scala 106:73]
  wire  _T_55 = _T_23 == 5'hb; // @[pe.scala 106:35]
  wire [4:0] _T_57 = _T_23 + 5'h1; // @[pe.scala 106:73]
  wire  _T_61 = _T_24 == 5'hb; // @[pe.scala 106:35]
  wire [4:0] _T_63 = _T_24 + 5'h1; // @[pe.scala 106:73]
  wire  _T_67 = _T_25 == 5'hb; // @[pe.scala 106:35]
  wire [4:0] _T_69 = _T_25 + 5'h1; // @[pe.scala 106:73]
  wire  _T_73 = _T_26 == 5'hb; // @[pe.scala 106:35]
  wire [4:0] _T_75 = _T_26 + 5'h1; // @[pe.scala 106:73]
  wire  _T_79 = _T_27 == 5'hb; // @[pe.scala 106:35]
  wire [4:0] _T_81 = _T_27 + 5'h1; // @[pe.scala 106:73]
  wire  _T_85 = _T_28 == 5'hb; // @[pe.scala 106:35]
  wire [4:0] _T_87 = _T_28 + 5'h1; // @[pe.scala 106:73]
  wire  _T_91 = _T_29 == 5'hb; // @[pe.scala 106:35]
  wire [4:0] _T_93 = _T_29 + 5'h1; // @[pe.scala 106:73]
  wire  _T_97 = _T_30 == 5'hb; // @[pe.scala 106:35]
  wire [4:0] _T_99 = _T_30 + 5'h1; // @[pe.scala 106:73]
  wire  _T_103 = _T_31 == 5'hb; // @[pe.scala 106:35]
  wire [4:0] _T_105 = _T_31 + 5'h1; // @[pe.scala 106:73]
  wire  _T_109 = _T_32 == 5'hb; // @[pe.scala 106:35]
  wire [4:0] _T_111 = _T_32 + 5'h1; // @[pe.scala 106:73]
  wire  _T_115 = _T_33 == 5'hb; // @[pe.scala 106:35]
  wire [4:0] _T_117 = _T_33 + 5'h1; // @[pe.scala 106:73]
  wire  _T_121 = _T_34 == 5'hb; // @[pe.scala 106:35]
  wire [4:0] _T_123 = _T_34 + 5'h1; // @[pe.scala 106:73]
  wire  _T_127 = _T_35 == 5'hb; // @[pe.scala 106:35]
  wire [4:0] _T_129 = _T_35 + 5'h1; // @[pe.scala 106:73]
  wire  _T_133 = _T_36 == 5'hb; // @[pe.scala 106:35]
  wire [4:0] _T_135 = _T_36 + 5'h1; // @[pe.scala 106:73]
  wire  _T_139 = _T_37 == 5'hb; // @[pe.scala 106:35]
  wire [4:0] _T_141 = _T_37 + 5'h1; // @[pe.scala 106:73]
  wire  _T_145 = _T_38 == 5'hb; // @[pe.scala 106:35]
  wire [4:0] _T_147 = _T_38 + 5'h1; // @[pe.scala 106:73]
  wire  _T_151 = _T_39 == 5'hb; // @[pe.scala 106:35]
  wire [4:0] _T_153 = _T_39 + 5'h1; // @[pe.scala 106:73]
  wire  _T_157 = _T_40 == 5'hb; // @[pe.scala 106:35]
  wire [4:0] _T_159 = _T_40 + 5'h1; // @[pe.scala 106:73]
  wire  _T_163 = _T_41 == 5'hb; // @[pe.scala 106:35]
  wire [4:0] _T_165 = _T_41 + 5'h1; // @[pe.scala 106:73]
  wire  _T_169 = _T_42 == 5'hb; // @[pe.scala 106:35]
  wire [4:0] _T_171 = _T_42 + 5'h1; // @[pe.scala 106:73]
  wire  _T_175 = _T_43 == 5'hb; // @[pe.scala 106:35]
  wire [4:0] _T_177 = _T_43 + 5'h1; // @[pe.scala 106:73]
  wire  _T_180 = _T_175 & io_to_pes_21_out_valid; // @[pe.scala 109:48]
  wire  _GEN_132 = _T_180 | _T_44; // @[pe.scala 109:81]
  wire  _T_181 = _T_45 == 10'hb; // @[pe.scala 113:29]
  wire [9:0] _T_183 = _T_45 + 10'h1; // @[pe.scala 113:65]
  wire  _T_186 = _T_46 == 10'h15; // @[pe.scala 114:61]
  wire [9:0] _T_188 = _T_46 + 10'h1; // @[pe.scala 114:94]
  wire  _T_193 = _T_181 & _T_186; // @[pe.scala 115:41]
  wire [127:0] _T_238_0 = _T__T_195_data; // @[pe.scala 119:32 pe.scala 119:32]
  wire [127:0] _T_238_1 = _T_1__T_197_data; // @[pe.scala 119:32 pe.scala 119:32]
  wire [127:0] _GEN_138 = 5'h1 == _T_46[4:0] ? _T_238_1 : _T_238_0; // @[pe.scala 121:20]
  wire [127:0] _T_238_2 = _T_2__T_199_data; // @[pe.scala 119:32 pe.scala 119:32]
  wire [127:0] _GEN_139 = 5'h2 == _T_46[4:0] ? _T_238_2 : _GEN_138; // @[pe.scala 121:20]
  wire [127:0] _T_238_3 = _T_3__T_201_data; // @[pe.scala 119:32 pe.scala 119:32]
  wire [127:0] _GEN_140 = 5'h3 == _T_46[4:0] ? _T_238_3 : _GEN_139; // @[pe.scala 121:20]
  wire [127:0] _T_238_4 = _T_4__T_203_data; // @[pe.scala 119:32 pe.scala 119:32]
  wire [127:0] _GEN_141 = 5'h4 == _T_46[4:0] ? _T_238_4 : _GEN_140; // @[pe.scala 121:20]
  wire [127:0] _T_238_5 = _T_5__T_205_data; // @[pe.scala 119:32 pe.scala 119:32]
  wire [127:0] _GEN_142 = 5'h5 == _T_46[4:0] ? _T_238_5 : _GEN_141; // @[pe.scala 121:20]
  wire [127:0] _T_238_6 = _T_6__T_207_data; // @[pe.scala 119:32 pe.scala 119:32]
  wire [127:0] _GEN_143 = 5'h6 == _T_46[4:0] ? _T_238_6 : _GEN_142; // @[pe.scala 121:20]
  wire [127:0] _T_238_7 = _T_7__T_209_data; // @[pe.scala 119:32 pe.scala 119:32]
  wire [127:0] _GEN_144 = 5'h7 == _T_46[4:0] ? _T_238_7 : _GEN_143; // @[pe.scala 121:20]
  wire [127:0] _T_238_8 = _T_8__T_211_data; // @[pe.scala 119:32 pe.scala 119:32]
  wire [127:0] _GEN_145 = 5'h8 == _T_46[4:0] ? _T_238_8 : _GEN_144; // @[pe.scala 121:20]
  wire [127:0] _T_238_9 = _T_9__T_213_data; // @[pe.scala 119:32 pe.scala 119:32]
  wire [127:0] _GEN_146 = 5'h9 == _T_46[4:0] ? _T_238_9 : _GEN_145; // @[pe.scala 121:20]
  wire [127:0] _T_238_10 = _T_10__T_215_data; // @[pe.scala 119:32 pe.scala 119:32]
  wire [127:0] _GEN_147 = 5'ha == _T_46[4:0] ? _T_238_10 : _GEN_146; // @[pe.scala 121:20]
  wire [127:0] _T_238_11 = _T_11__T_217_data; // @[pe.scala 119:32 pe.scala 119:32]
  wire [127:0] _GEN_148 = 5'hb == _T_46[4:0] ? _T_238_11 : _GEN_147; // @[pe.scala 121:20]
  wire [127:0] _T_238_12 = _T_12__T_219_data; // @[pe.scala 119:32 pe.scala 119:32]
  wire [127:0] _GEN_149 = 5'hc == _T_46[4:0] ? _T_238_12 : _GEN_148; // @[pe.scala 121:20]
  wire [127:0] _T_238_13 = _T_13__T_221_data; // @[pe.scala 119:32 pe.scala 119:32]
  wire [127:0] _GEN_150 = 5'hd == _T_46[4:0] ? _T_238_13 : _GEN_149; // @[pe.scala 121:20]
  wire [127:0] _T_238_14 = _T_14__T_223_data; // @[pe.scala 119:32 pe.scala 119:32]
  wire [127:0] _GEN_151 = 5'he == _T_46[4:0] ? _T_238_14 : _GEN_150; // @[pe.scala 121:20]
  wire [127:0] _T_238_15 = _T_15__T_225_data; // @[pe.scala 119:32 pe.scala 119:32]
  wire [127:0] _GEN_152 = 5'hf == _T_46[4:0] ? _T_238_15 : _GEN_151; // @[pe.scala 121:20]
  wire [127:0] _T_238_16 = _T_16__T_227_data; // @[pe.scala 119:32 pe.scala 119:32]
  wire [127:0] _GEN_153 = 5'h10 == _T_46[4:0] ? _T_238_16 : _GEN_152; // @[pe.scala 121:20]
  wire [127:0] _T_238_17 = _T_17__T_229_data; // @[pe.scala 119:32 pe.scala 119:32]
  wire [127:0] _GEN_154 = 5'h11 == _T_46[4:0] ? _T_238_17 : _GEN_153; // @[pe.scala 121:20]
  wire [127:0] _T_238_18 = _T_18__T_231_data; // @[pe.scala 119:32 pe.scala 119:32]
  wire [127:0] _GEN_155 = 5'h12 == _T_46[4:0] ? _T_238_18 : _GEN_154; // @[pe.scala 121:20]
  wire [127:0] _T_238_19 = _T_19__T_233_data; // @[pe.scala 119:32 pe.scala 119:32]
  wire [127:0] _GEN_156 = 5'h13 == _T_46[4:0] ? _T_238_19 : _GEN_155; // @[pe.scala 121:20]
  wire [127:0] _T_238_20 = _T_20__T_235_data; // @[pe.scala 119:32 pe.scala 119:32]
  wire [127:0] _GEN_157 = 5'h14 == _T_46[4:0] ? _T_238_20 : _GEN_156; // @[pe.scala 121:20]
  wire [127:0] _T_238_21 = _T_21__T_237_data; // @[pe.scala 119:32 pe.scala 119:32]
  reg  _T_240; // @[Reg.scala 15:16]
  reg [31:0] _RAND_113;
  reg  _T_241; // @[Reg.scala 15:16]
  reg [31:0] _RAND_114;
  reg  _T_242; // @[Reg.scala 15:16]
  reg [31:0] _RAND_115;
  reg  _T_243; // @[Reg.scala 15:16]
  reg [31:0] _RAND_116;
  reg  _T_244; // @[Reg.scala 15:16]
  reg [31:0] _RAND_117;
  reg  _T_245; // @[Reg.scala 15:16]
  reg [31:0] _RAND_118;
  reg  _T_246; // @[Reg.scala 15:16]
  reg [31:0] _RAND_119;
  reg  _T_247; // @[Reg.scala 15:16]
  reg [31:0] _RAND_120;
  reg  _T_248; // @[Reg.scala 15:16]
  reg [31:0] _RAND_121;
  reg  _T_249; // @[Reg.scala 15:16]
  reg [31:0] _RAND_122;
  reg  _T_250; // @[Reg.scala 15:16]
  reg [31:0] _RAND_123;
  reg  _T_251; // @[Reg.scala 15:16]
  reg [31:0] _RAND_124;
  reg  _T_252; // @[Reg.scala 15:16]
  reg [31:0] _RAND_125;
  reg  _T_253; // @[Reg.scala 15:16]
  reg [31:0] _RAND_126;
  reg  _T_254; // @[Reg.scala 15:16]
  reg [31:0] _RAND_127;
  reg  _T_255; // @[Reg.scala 15:16]
  reg [31:0] _RAND_128;
  reg  _T_256; // @[Reg.scala 15:16]
  reg [31:0] _RAND_129;
  reg  _T_257; // @[Reg.scala 15:16]
  reg [31:0] _RAND_130;
  reg  _T_258; // @[Reg.scala 15:16]
  reg [31:0] _RAND_131;
  reg  _T_259; // @[Reg.scala 15:16]
  reg [31:0] _RAND_132;
  reg  _T_260; // @[Reg.scala 15:16]
  reg [31:0] _RAND_133;
  reg  _T_261; // @[Reg.scala 15:16]
  reg [31:0] _RAND_134;
  reg  _T_262; // @[Reg.scala 15:16]
  reg [31:0] _RAND_135;
  reg  _T_263; // @[Reg.scala 15:16]
  reg [31:0] _RAND_136;
  reg  _T_264; // @[Reg.scala 15:16]
  reg [31:0] _RAND_137;
  reg  _T_265; // @[Reg.scala 15:16]
  reg [31:0] _RAND_138;
  reg  _T_266; // @[Reg.scala 15:16]
  reg [31:0] _RAND_139;
  reg  _T_267; // @[Reg.scala 15:16]
  reg [31:0] _RAND_140;
  reg  _T_268; // @[Reg.scala 15:16]
  reg [31:0] _RAND_141;
  reg  _T_269; // @[Reg.scala 15:16]
  reg [31:0] _RAND_142;
  reg  _T_270; // @[Reg.scala 15:16]
  reg [31:0] _RAND_143;
  reg  _T_271; // @[Reg.scala 15:16]
  reg [31:0] _RAND_144;
  reg  _T_272; // @[Reg.scala 15:16]
  reg [31:0] _RAND_145;
  reg  _T_273; // @[Reg.scala 15:16]
  reg [31:0] _RAND_146;
  reg  _T_274; // @[Reg.scala 15:16]
  reg [31:0] _RAND_147;
  reg  _T_275; // @[Reg.scala 15:16]
  reg [31:0] _RAND_148;
  reg  _T_276; // @[Reg.scala 15:16]
  reg [31:0] _RAND_149;
  reg  _T_277; // @[Reg.scala 15:16]
  reg [31:0] _RAND_150;
  reg  _T_278; // @[Reg.scala 15:16]
  reg [31:0] _RAND_151;
  reg  _T_279; // @[Reg.scala 15:16]
  reg [31:0] _RAND_152;
  reg  _T_280; // @[Reg.scala 15:16]
  reg [31:0] _RAND_153;
  reg  _T_281; // @[Reg.scala 15:16]
  reg [31:0] _RAND_154;
  reg  _T_282; // @[Reg.scala 15:16]
  reg [31:0] _RAND_155;
  reg  _T_283; // @[Reg.scala 15:16]
  reg [31:0] _RAND_156;
  reg  _T_284; // @[Reg.scala 15:16]
  reg [31:0] _RAND_157;
  reg  _T_285; // @[Reg.scala 15:16]
  reg [31:0] _RAND_158;
  reg  _T_286; // @[Reg.scala 15:16]
  reg [31:0] _RAND_159;
  reg  _T_287; // @[Reg.scala 15:16]
  reg [31:0] _RAND_160;
  reg  _T_288; // @[Reg.scala 15:16]
  reg [31:0] _RAND_161;
  reg  _T_289; // @[Reg.scala 15:16]
  reg [31:0] _RAND_162;
  reg  _T_290; // @[Reg.scala 15:16]
  reg [31:0] _RAND_163;
  reg  _T_291; // @[Reg.scala 15:16]
  reg [31:0] _RAND_164;
  reg  _T_292; // @[Reg.scala 15:16]
  reg [31:0] _RAND_165;
  reg  _T_293; // @[Reg.scala 15:16]
  reg [31:0] _RAND_166;
  reg  _T_294; // @[Reg.scala 15:16]
  reg [31:0] _RAND_167;
  reg  _T_295; // @[Reg.scala 15:16]
  reg [31:0] _RAND_168;
  reg  _T_296; // @[Reg.scala 15:16]
  reg [31:0] _RAND_169;
  reg  _T_297; // @[Reg.scala 15:16]
  reg [31:0] _RAND_170;
  reg  _T_298; // @[Reg.scala 15:16]
  reg [31:0] _RAND_171;
  reg  _T_299; // @[Reg.scala 15:16]
  reg [31:0] _RAND_172;
  reg  _T_300; // @[Reg.scala 15:16]
  reg [31:0] _RAND_173;
  reg  _T_301; // @[Reg.scala 15:16]
  reg [31:0] _RAND_174;
  reg  _T_302; // @[Reg.scala 15:16]
  reg [31:0] _RAND_175;
  reg  _T_303; // @[Reg.scala 15:16]
  reg [31:0] _RAND_176;
  reg  _T_304; // @[Reg.scala 15:16]
  reg [31:0] _RAND_177;
  reg  _T_305; // @[Reg.scala 15:16]
  reg [31:0] _RAND_178;
  reg  _T_306; // @[Reg.scala 15:16]
  reg [31:0] _RAND_179;
  reg  _T_307; // @[Reg.scala 15:16]
  reg [31:0] _RAND_180;
  reg  _T_308; // @[Reg.scala 15:16]
  reg [31:0] _RAND_181;
  reg  _T_309; // @[Reg.scala 15:16]
  reg [31:0] _RAND_182;
  reg  _T_310; // @[Reg.scala 15:16]
  reg [31:0] _RAND_183;
  reg  _T_311; // @[Reg.scala 15:16]
  reg [31:0] _RAND_184;
  reg  _T_312; // @[Reg.scala 15:16]
  reg [31:0] _RAND_185;
  reg  _T_313; // @[Reg.scala 15:16]
  reg [31:0] _RAND_186;
  reg  _T_314; // @[Reg.scala 15:16]
  reg [31:0] _RAND_187;
  reg  _T_315; // @[Reg.scala 15:16]
  reg [31:0] _RAND_188;
  reg  _T_316; // @[Reg.scala 15:16]
  reg [31:0] _RAND_189;
  reg  _T_317; // @[Reg.scala 15:16]
  reg [31:0] _RAND_190;
  reg  _T_318; // @[Reg.scala 15:16]
  reg [31:0] _RAND_191;
  reg  _T_319; // @[Reg.scala 15:16]
  reg [31:0] _RAND_192;
  reg  _T_320; // @[Reg.scala 15:16]
  reg [31:0] _RAND_193;
  reg  _T_321; // @[Reg.scala 15:16]
  reg [31:0] _RAND_194;
  reg  _T_322; // @[Reg.scala 15:16]
  reg [31:0] _RAND_195;
  reg  _T_323; // @[Reg.scala 15:16]
  reg [31:0] _RAND_196;
  reg  _T_324; // @[Reg.scala 15:16]
  reg [31:0] _RAND_197;
  reg  _T_325; // @[Reg.scala 15:16]
  reg [31:0] _RAND_198;
  reg  _T_326; // @[Reg.scala 15:16]
  reg [31:0] _RAND_199;
  reg  _T_327; // @[Reg.scala 15:16]
  reg [31:0] _RAND_200;
  reg  _T_328; // @[Reg.scala 15:16]
  reg [31:0] _RAND_201;
  reg  _T_329; // @[Reg.scala 15:16]
  reg [31:0] _RAND_202;
  reg  _T_330; // @[Reg.scala 15:16]
  reg [31:0] _RAND_203;
  reg  _T_331; // @[Reg.scala 15:16]
  reg [31:0] _RAND_204;
  reg  _T_332; // @[Reg.scala 15:16]
  reg [31:0] _RAND_205;
  reg  _T_333; // @[Reg.scala 15:16]
  reg [31:0] _RAND_206;
  reg  _T_334; // @[Reg.scala 15:16]
  reg [31:0] _RAND_207;
  reg  _T_335; // @[Reg.scala 15:16]
  reg [31:0] _RAND_208;
  reg  _T_336; // @[Reg.scala 15:16]
  reg [31:0] _RAND_209;
  reg  _T_337; // @[Reg.scala 15:16]
  reg [31:0] _RAND_210;
  reg  _T_338; // @[Reg.scala 15:16]
  reg [31:0] _RAND_211;
  reg  _T_339; // @[Reg.scala 15:16]
  reg [31:0] _RAND_212;
  reg  _T_340; // @[Reg.scala 15:16]
  reg [31:0] _RAND_213;
  reg  _T_341; // @[Reg.scala 15:16]
  reg [31:0] _RAND_214;
  reg  _T_342; // @[Reg.scala 15:16]
  reg [31:0] _RAND_215;
  reg  _T_343; // @[Reg.scala 15:16]
  reg [31:0] _RAND_216;
  reg  _T_344; // @[Reg.scala 15:16]
  reg [31:0] _RAND_217;
  reg  _T_345; // @[Reg.scala 15:16]
  reg [31:0] _RAND_218;
  reg  _T_346; // @[Reg.scala 15:16]
  reg [31:0] _RAND_219;
  reg  _T_347; // @[Reg.scala 15:16]
  reg [31:0] _RAND_220;
  reg  _T_348; // @[Reg.scala 15:16]
  reg [31:0] _RAND_221;
  reg  _T_349; // @[Reg.scala 15:16]
  reg [31:0] _RAND_222;
  reg  _T_350; // @[Reg.scala 15:16]
  reg [31:0] _RAND_223;
  reg  _T_351; // @[Reg.scala 15:16]
  reg [31:0] _RAND_224;
  reg  _T_352; // @[Reg.scala 15:16]
  reg [31:0] _RAND_225;
  reg  _T_353; // @[Reg.scala 15:16]
  reg [31:0] _RAND_226;
  reg  _T_354; // @[Reg.scala 15:16]
  reg [31:0] _RAND_227;
  reg  _T_355; // @[Reg.scala 15:16]
  reg [31:0] _RAND_228;
  reg  _T_356; // @[Reg.scala 15:16]
  reg [31:0] _RAND_229;
  reg  _T_357; // @[Reg.scala 15:16]
  reg [31:0] _RAND_230;
  reg  _T_358; // @[Reg.scala 15:16]
  reg [31:0] _RAND_231;
  reg  _T_359; // @[Reg.scala 15:16]
  reg [31:0] _RAND_232;
  reg  _T_360; // @[Reg.scala 15:16]
  reg [31:0] _RAND_233;
  reg  _T_361; // @[Reg.scala 15:16]
  reg [31:0] _RAND_234;
  reg  _T_362; // @[Reg.scala 15:16]
  reg [31:0] _RAND_235;
  reg  _T_363; // @[Reg.scala 15:16]
  reg [31:0] _RAND_236;
  reg  _T_364; // @[Reg.scala 15:16]
  reg [31:0] _RAND_237;
  reg  _T_365; // @[Reg.scala 15:16]
  reg [31:0] _RAND_238;
  reg  _T_366; // @[Reg.scala 15:16]
  reg [31:0] _RAND_239;
  reg  _T_367; // @[Reg.scala 15:16]
  reg [31:0] _RAND_240;
  reg  _T_368; // @[Reg.scala 15:16]
  reg [31:0] _RAND_241;
  reg  _T_369; // @[Reg.scala 15:16]
  reg [31:0] _RAND_242;
  reg  _T_370; // @[Reg.scala 15:16]
  reg [31:0] _RAND_243;
  reg  _T_371; // @[Reg.scala 15:16]
  reg [31:0] _RAND_244;
  reg  _T_372; // @[Reg.scala 15:16]
  reg [31:0] _RAND_245;
  reg  _T_373; // @[Reg.scala 15:16]
  reg [31:0] _RAND_246;
  reg  _T_374; // @[Reg.scala 15:16]
  reg [31:0] _RAND_247;
  reg  _T_375; // @[Reg.scala 15:16]
  reg [31:0] _RAND_248;
  reg  _T_376; // @[Reg.scala 15:16]
  reg [31:0] _RAND_249;
  reg  _T_377; // @[Reg.scala 15:16]
  reg [31:0] _RAND_250;
  reg  _T_378; // @[Reg.scala 15:16]
  reg [31:0] _RAND_251;
  reg  _T_379; // @[Reg.scala 15:16]
  reg [31:0] _RAND_252;
  reg  _T_380; // @[Reg.scala 15:16]
  reg [31:0] _RAND_253;
  reg  _T_381; // @[Reg.scala 15:16]
  reg [31:0] _RAND_254;
  reg  _T_382; // @[Reg.scala 15:16]
  reg [31:0] _RAND_255;
  reg  _T_383; // @[Reg.scala 15:16]
  reg [31:0] _RAND_256;
  reg  _T_384; // @[Reg.scala 15:16]
  reg [31:0] _RAND_257;
  reg  _T_385; // @[Reg.scala 15:16]
  reg [31:0] _RAND_258;
  reg  _T_386; // @[Reg.scala 15:16]
  reg [31:0] _RAND_259;
  reg  _T_387; // @[Reg.scala 15:16]
  reg [31:0] _RAND_260;
  reg  _T_388; // @[Reg.scala 15:16]
  reg [31:0] _RAND_261;
  reg  _T_389; // @[Reg.scala 15:16]
  reg [31:0] _RAND_262;
  reg  _T_390; // @[Reg.scala 15:16]
  reg [31:0] _RAND_263;
  reg  _T_391; // @[Reg.scala 15:16]
  reg [31:0] _RAND_264;
  reg  _T_392; // @[Reg.scala 15:16]
  reg [31:0] _RAND_265;
  reg  _T_393; // @[Reg.scala 15:16]
  reg [31:0] _RAND_266;
  reg  _T_394; // @[Reg.scala 15:16]
  reg [31:0] _RAND_267;
  reg  _T_395; // @[Reg.scala 15:16]
  reg [31:0] _RAND_268;
  reg  _T_396; // @[Reg.scala 15:16]
  reg [31:0] _RAND_269;
  reg  _T_397; // @[Reg.scala 15:16]
  reg [31:0] _RAND_270;
  reg  _T_398; // @[Reg.scala 15:16]
  reg [31:0] _RAND_271;
  reg  _T_399; // @[Reg.scala 15:16]
  reg [31:0] _RAND_272;
  reg  _T_400; // @[Reg.scala 15:16]
  reg [31:0] _RAND_273;
  reg  _T_401; // @[Reg.scala 15:16]
  reg [31:0] _RAND_274;
  reg  _T_402; // @[Reg.scala 15:16]
  reg [31:0] _RAND_275;
  reg  _T_403; // @[Reg.scala 15:16]
  reg [31:0] _RAND_276;
  reg  _T_404; // @[Reg.scala 15:16]
  reg [31:0] _RAND_277;
  reg  _T_405; // @[Reg.scala 15:16]
  reg [31:0] _RAND_278;
  reg  _T_406; // @[Reg.scala 15:16]
  reg [31:0] _RAND_279;
  reg  _T_407; // @[Reg.scala 15:16]
  reg [31:0] _RAND_280;
  reg  _T_408; // @[Reg.scala 15:16]
  reg [31:0] _RAND_281;
  reg  _T_409; // @[Reg.scala 15:16]
  reg [31:0] _RAND_282;
  reg  _T_410; // @[Reg.scala 15:16]
  reg [31:0] _RAND_283;
  reg  _T_411; // @[Reg.scala 15:16]
  reg [31:0] _RAND_284;
  reg  _T_412; // @[Reg.scala 15:16]
  reg [31:0] _RAND_285;
  reg  _T_413; // @[Reg.scala 15:16]
  reg [31:0] _RAND_286;
  reg  _T_414; // @[Reg.scala 15:16]
  reg [31:0] _RAND_287;
  reg  _T_415; // @[Reg.scala 15:16]
  reg [31:0] _RAND_288;
  reg  _T_416; // @[Reg.scala 15:16]
  reg [31:0] _RAND_289;
  reg  _T_417; // @[Reg.scala 15:16]
  reg [31:0] _RAND_290;
  reg  _T_418; // @[Reg.scala 15:16]
  reg [31:0] _RAND_291;
  reg  _T_419; // @[Reg.scala 15:16]
  reg [31:0] _RAND_292;
  reg  _T_420; // @[Reg.scala 15:16]
  reg [31:0] _RAND_293;
  reg  _T_421; // @[Reg.scala 15:16]
  reg [31:0] _RAND_294;
  reg  _T_422; // @[Reg.scala 15:16]
  reg [31:0] _RAND_295;
  reg  _T_423; // @[Reg.scala 15:16]
  reg [31:0] _RAND_296;
  reg  _T_424; // @[Reg.scala 15:16]
  reg [31:0] _RAND_297;
  reg  _T_425; // @[Reg.scala 15:16]
  reg [31:0] _RAND_298;
  reg  _T_426; // @[Reg.scala 15:16]
  reg [31:0] _RAND_299;
  reg  _T_427; // @[Reg.scala 15:16]
  reg [31:0] _RAND_300;
  reg  _T_428; // @[Reg.scala 15:16]
  reg [31:0] _RAND_301;
  reg  _T_429; // @[Reg.scala 15:16]
  reg [31:0] _RAND_302;
  reg  _T_430; // @[Reg.scala 15:16]
  reg [31:0] _RAND_303;
  reg  _T_431; // @[Reg.scala 15:16]
  reg [31:0] _RAND_304;
  reg  _T_432; // @[Reg.scala 15:16]
  reg [31:0] _RAND_305;
  reg  _T_433; // @[Reg.scala 15:16]
  reg [31:0] _RAND_306;
  reg  _T_434; // @[Reg.scala 15:16]
  reg [31:0] _RAND_307;
  reg  _T_435; // @[Reg.scala 15:16]
  reg [31:0] _RAND_308;
  reg  _T_436; // @[Reg.scala 15:16]
  reg [31:0] _RAND_309;
  reg  _T_437; // @[Reg.scala 15:16]
  reg [31:0] _RAND_310;
  reg  _T_438; // @[Reg.scala 15:16]
  reg [31:0] _RAND_311;
  reg  _T_439; // @[Reg.scala 15:16]
  reg [31:0] _RAND_312;
  reg  _T_440; // @[Reg.scala 15:16]
  reg [31:0] _RAND_313;
  reg  _T_441; // @[Reg.scala 15:16]
  reg [31:0] _RAND_314;
  reg  _T_442; // @[Reg.scala 15:16]
  reg [31:0] _RAND_315;
  reg  _T_443; // @[Reg.scala 15:16]
  reg [31:0] _RAND_316;
  reg  _T_444; // @[Reg.scala 15:16]
  reg [31:0] _RAND_317;
  reg  _T_445; // @[Reg.scala 15:16]
  reg [31:0] _RAND_318;
  reg  _T_446; // @[Reg.scala 15:16]
  reg [31:0] _RAND_319;
  reg  _T_447; // @[Reg.scala 15:16]
  reg [31:0] _RAND_320;
  reg  _T_448; // @[Reg.scala 15:16]
  reg [31:0] _RAND_321;
  reg  _T_449; // @[Reg.scala 15:16]
  reg [31:0] _RAND_322;
  reg  _T_450; // @[Reg.scala 15:16]
  reg [31:0] _RAND_323;
  reg  _T_451; // @[Reg.scala 15:16]
  reg [31:0] _RAND_324;
  reg  _T_452; // @[Reg.scala 15:16]
  reg [31:0] _RAND_325;
  reg  _T_453; // @[Reg.scala 15:16]
  reg [31:0] _RAND_326;
  reg  _T_454; // @[Reg.scala 15:16]
  reg [31:0] _RAND_327;
  reg  _T_455; // @[Reg.scala 15:16]
  reg [31:0] _RAND_328;
  reg  _T_456; // @[Reg.scala 15:16]
  reg [31:0] _RAND_329;
  reg  _T_457; // @[Reg.scala 15:16]
  reg [31:0] _RAND_330;
  reg  _T_458; // @[Reg.scala 15:16]
  reg [31:0] _RAND_331;
  reg  _T_459; // @[Reg.scala 15:16]
  reg [31:0] _RAND_332;
  reg  _T_460; // @[Reg.scala 15:16]
  reg [31:0] _RAND_333;
  reg  _T_461; // @[Reg.scala 15:16]
  reg [31:0] _RAND_334;
  reg  _T_462; // @[Reg.scala 15:16]
  reg [31:0] _RAND_335;
  reg  _T_463; // @[Reg.scala 15:16]
  reg [31:0] _RAND_336;
  reg  _T_464; // @[Reg.scala 15:16]
  reg [31:0] _RAND_337;
  reg  _T_465; // @[Reg.scala 15:16]
  reg [31:0] _RAND_338;
  reg  _T_466; // @[Reg.scala 15:16]
  reg [31:0] _RAND_339;
  reg  _T_467; // @[Reg.scala 15:16]
  reg [31:0] _RAND_340;
  reg  _T_468; // @[Reg.scala 15:16]
  reg [31:0] _RAND_341;
  reg  _T_469; // @[Reg.scala 15:16]
  reg [31:0] _RAND_342;
  reg  _T_470; // @[Reg.scala 15:16]
  reg [31:0] _RAND_343;
  reg  _T_471; // @[Reg.scala 15:16]
  reg [31:0] _RAND_344;
  reg  _T_472; // @[Reg.scala 15:16]
  reg [31:0] _RAND_345;
  reg  _T_473; // @[Reg.scala 15:16]
  reg [31:0] _RAND_346;
  reg  _T_474; // @[Reg.scala 15:16]
  reg [31:0] _RAND_347;
  reg  _T_475; // @[Reg.scala 15:16]
  reg [31:0] _RAND_348;
  reg  _T_476; // @[Reg.scala 15:16]
  reg [31:0] _RAND_349;
  reg  _T_477; // @[Reg.scala 15:16]
  reg [31:0] _RAND_350;
  reg  _T_478; // @[Reg.scala 15:16]
  reg [31:0] _RAND_351;
  reg  _T_479; // @[Reg.scala 15:16]
  reg [31:0] _RAND_352;
  reg  _T_480; // @[Reg.scala 15:16]
  reg [31:0] _RAND_353;
  reg  _T_481; // @[Reg.scala 15:16]
  reg [31:0] _RAND_354;
  reg  _T_482; // @[Reg.scala 15:16]
  reg [31:0] _RAND_355;
  reg  _T_483; // @[Reg.scala 15:16]
  reg [31:0] _RAND_356;
  reg  _T_484; // @[Reg.scala 15:16]
  reg [31:0] _RAND_357;
  reg  _T_485; // @[Reg.scala 15:16]
  reg [31:0] _RAND_358;
  reg  _T_486; // @[Reg.scala 15:16]
  reg [31:0] _RAND_359;
  reg  _T_487; // @[Reg.scala 15:16]
  reg [31:0] _RAND_360;
  reg  _T_488; // @[Reg.scala 15:16]
  reg [31:0] _RAND_361;
  reg  _T_489; // @[Reg.scala 15:16]
  reg [31:0] _RAND_362;
  reg  _T_490; // @[Reg.scala 15:16]
  reg [31:0] _RAND_363;
  reg  _T_491; // @[Reg.scala 15:16]
  reg [31:0] _RAND_364;
  reg  _T_492; // @[Reg.scala 15:16]
  reg [31:0] _RAND_365;
  reg  _T_493; // @[Reg.scala 15:16]
  reg [31:0] _RAND_366;
  reg  _T_494; // @[Reg.scala 15:16]
  reg [31:0] _RAND_367;
  reg  _T_495; // @[Reg.scala 15:16]
  reg [31:0] _RAND_368;
  reg  _T_496; // @[Reg.scala 15:16]
  reg [31:0] _RAND_369;
  reg  _T_497; // @[Reg.scala 15:16]
  reg [31:0] _RAND_370;
  reg  _T_498; // @[Reg.scala 15:16]
  reg [31:0] _RAND_371;
  reg  _T_499; // @[Reg.scala 15:16]
  reg [31:0] _RAND_372;
  reg  _T_500; // @[Reg.scala 15:16]
  reg [31:0] _RAND_373;
  reg  _T_501; // @[Reg.scala 15:16]
  reg [31:0] _RAND_374;
  reg  _T_502; // @[Reg.scala 15:16]
  reg [31:0] _RAND_375;
  reg  _T_503; // @[Reg.scala 15:16]
  reg [31:0] _RAND_376;
  reg  _T_504; // @[Reg.scala 15:16]
  reg [31:0] _RAND_377;
  reg  _T_505; // @[Reg.scala 15:16]
  reg [31:0] _RAND_378;
  reg  _T_506; // @[Reg.scala 15:16]
  reg [31:0] _RAND_379;
  reg  _T_507; // @[Reg.scala 15:16]
  reg [31:0] _RAND_380;
  reg  _T_508; // @[Reg.scala 15:16]
  reg [31:0] _RAND_381;
  reg  _T_509; // @[Reg.scala 15:16]
  reg [31:0] _RAND_382;
  reg  _T_510; // @[Reg.scala 15:16]
  reg [31:0] _RAND_383;
  reg  _T_511; // @[Reg.scala 15:16]
  reg [31:0] _RAND_384;
  reg  _T_512; // @[Reg.scala 15:16]
  reg [31:0] _RAND_385;
  reg  _T_513; // @[Reg.scala 15:16]
  reg [31:0] _RAND_386;
  reg  _T_514; // @[Reg.scala 15:16]
  reg [31:0] _RAND_387;
  reg  _T_515; // @[Reg.scala 15:16]
  reg [31:0] _RAND_388;
  reg  _T_516; // @[Reg.scala 15:16]
  reg [31:0] _RAND_389;
  reg  _T_517; // @[Reg.scala 15:16]
  reg [31:0] _RAND_390;
  reg  _T_518; // @[Reg.scala 15:16]
  reg [31:0] _RAND_391;
  reg  _T_519; // @[Reg.scala 15:16]
  reg [31:0] _RAND_392;
  reg  _T_520; // @[Reg.scala 15:16]
  reg [31:0] _RAND_393;
  reg  _T_521; // @[Reg.scala 15:16]
  reg [31:0] _RAND_394;
  reg  _T_522; // @[Reg.scala 15:16]
  reg [31:0] _RAND_395;
  reg  _T_523; // @[Reg.scala 15:16]
  reg [31:0] _RAND_396;
  reg  _T_524; // @[Reg.scala 15:16]
  reg [31:0] _RAND_397;
  reg  _T_525; // @[Reg.scala 15:16]
  reg [31:0] _RAND_398;
  reg  _T_526; // @[Reg.scala 15:16]
  reg [31:0] _RAND_399;
  reg  _T_527; // @[Reg.scala 15:16]
  reg [31:0] _RAND_400;
  reg  _T_528; // @[Reg.scala 15:16]
  reg [31:0] _RAND_401;
  reg  _T_529; // @[Reg.scala 15:16]
  reg [31:0] _RAND_402;
  reg  _T_530; // @[Reg.scala 15:16]
  reg [31:0] _RAND_403;
  reg  _T_531; // @[Reg.scala 15:16]
  reg [31:0] _RAND_404;
  reg  _T_532; // @[Reg.scala 15:16]
  reg [31:0] _RAND_405;
  reg  _T_533; // @[Reg.scala 15:16]
  reg [31:0] _RAND_406;
  reg  _T_534; // @[Reg.scala 15:16]
  reg [31:0] _RAND_407;
  reg  _T_535; // @[Reg.scala 15:16]
  reg [31:0] _RAND_408;
  reg  _T_536; // @[Reg.scala 15:16]
  reg [31:0] _RAND_409;
  reg  _T_537; // @[Reg.scala 15:16]
  reg [31:0] _RAND_410;
  reg  _T_538; // @[Reg.scala 15:16]
  reg [31:0] _RAND_411;
  reg  _T_539; // @[Reg.scala 15:16]
  reg [31:0] _RAND_412;
  reg  _T_540; // @[Reg.scala 15:16]
  reg [31:0] _RAND_413;
  reg  _T_541; // @[Reg.scala 15:16]
  reg [31:0] _RAND_414;
  reg  _T_542; // @[Reg.scala 15:16]
  reg [31:0] _RAND_415;
  reg  _T_543; // @[Reg.scala 15:16]
  reg [31:0] _RAND_416;
  reg  _T_544; // @[Reg.scala 15:16]
  reg [31:0] _RAND_417;
  reg  _T_545; // @[Reg.scala 15:16]
  reg [31:0] _RAND_418;
  reg  _T_546; // @[Reg.scala 15:16]
  reg [31:0] _RAND_419;
  reg  _T_547; // @[Reg.scala 15:16]
  reg [31:0] _RAND_420;
  reg  _T_548; // @[Reg.scala 15:16]
  reg [31:0] _RAND_421;
  reg  _T_549; // @[Reg.scala 15:16]
  reg [31:0] _RAND_422;
  reg  _T_550; // @[Reg.scala 15:16]
  reg [31:0] _RAND_423;
  reg  _T_551; // @[Reg.scala 15:16]
  reg [31:0] _RAND_424;
  reg  _T_552; // @[Reg.scala 15:16]
  reg [31:0] _RAND_425;
  reg  _T_553; // @[Reg.scala 15:16]
  reg [31:0] _RAND_426;
  reg  _T_554; // @[Reg.scala 15:16]
  reg [31:0] _RAND_427;
  reg  _T_555; // @[Reg.scala 15:16]
  reg [31:0] _RAND_428;
  reg  _T_556; // @[Reg.scala 15:16]
  reg [31:0] _RAND_429;
  reg  _T_557; // @[Reg.scala 15:16]
  reg [31:0] _RAND_430;
  reg  _T_558; // @[Reg.scala 15:16]
  reg [31:0] _RAND_431;
  reg  _T_559; // @[Reg.scala 15:16]
  reg [31:0] _RAND_432;
  reg  _T_560; // @[Reg.scala 15:16]
  reg [31:0] _RAND_433;
  reg  _T_561; // @[Reg.scala 15:16]
  reg [31:0] _RAND_434;
  reg  _T_562; // @[Reg.scala 15:16]
  reg [31:0] _RAND_435;
  reg  _T_563; // @[Reg.scala 15:16]
  reg [31:0] _RAND_436;
  reg  _T_564; // @[Reg.scala 15:16]
  reg [31:0] _RAND_437;
  reg  _T_565; // @[Reg.scala 15:16]
  reg [31:0] _RAND_438;
  reg  _T_566; // @[Reg.scala 15:16]
  reg [31:0] _RAND_439;
  reg  _T_567; // @[Reg.scala 15:16]
  reg [31:0] _RAND_440;
  reg  _T_568; // @[Reg.scala 15:16]
  reg [31:0] _RAND_441;
  reg  _T_569; // @[Reg.scala 15:16]
  reg [31:0] _RAND_442;
  assign _T__T_195_addr = _T__T_195_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T__T_195_data = _T[_T__T_195_addr]; // @[pe.scala 94:49]
  `else
  assign _T__T_195_data = _T__T_195_addr >= 4'hc ? _RAND_1[127:0] : _T[_T__T_195_addr]; // @[pe.scala 94:49]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T__T_48_data = io_to_pes_0_out_bits;
  assign _T__T_48_addr = _T_22[3:0];
  assign _T__T_48_mask = 1'h1;
  assign _T__T_48_en = io_to_pes_0_out_valid;
  assign _T_1__T_197_addr = _T_1__T_197_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_1__T_197_data = _T_1[_T_1__T_197_addr]; // @[pe.scala 94:49]
  `else
  assign _T_1__T_197_data = _T_1__T_197_addr >= 4'hc ? _RAND_5[127:0] : _T_1[_T_1__T_197_addr]; // @[pe.scala 94:49]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_1__T_54_data = io_to_pes_1_out_bits;
  assign _T_1__T_54_addr = _T_23[3:0];
  assign _T_1__T_54_mask = 1'h1;
  assign _T_1__T_54_en = io_to_pes_1_out_valid;
  assign _T_2__T_199_addr = _T_2__T_199_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_2__T_199_data = _T_2[_T_2__T_199_addr]; // @[pe.scala 94:49]
  `else
  assign _T_2__T_199_data = _T_2__T_199_addr >= 4'hc ? _RAND_9[127:0] : _T_2[_T_2__T_199_addr]; // @[pe.scala 94:49]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_2__T_60_data = io_to_pes_2_out_bits;
  assign _T_2__T_60_addr = _T_24[3:0];
  assign _T_2__T_60_mask = 1'h1;
  assign _T_2__T_60_en = io_to_pes_2_out_valid;
  assign _T_3__T_201_addr = _T_3__T_201_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_3__T_201_data = _T_3[_T_3__T_201_addr]; // @[pe.scala 94:49]
  `else
  assign _T_3__T_201_data = _T_3__T_201_addr >= 4'hc ? _RAND_13[127:0] : _T_3[_T_3__T_201_addr]; // @[pe.scala 94:49]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_3__T_66_data = io_to_pes_3_out_bits;
  assign _T_3__T_66_addr = _T_25[3:0];
  assign _T_3__T_66_mask = 1'h1;
  assign _T_3__T_66_en = io_to_pes_3_out_valid;
  assign _T_4__T_203_addr = _T_4__T_203_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_4__T_203_data = _T_4[_T_4__T_203_addr]; // @[pe.scala 94:49]
  `else
  assign _T_4__T_203_data = _T_4__T_203_addr >= 4'hc ? _RAND_17[127:0] : _T_4[_T_4__T_203_addr]; // @[pe.scala 94:49]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_4__T_72_data = io_to_pes_4_out_bits;
  assign _T_4__T_72_addr = _T_26[3:0];
  assign _T_4__T_72_mask = 1'h1;
  assign _T_4__T_72_en = io_to_pes_4_out_valid;
  assign _T_5__T_205_addr = _T_5__T_205_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_5__T_205_data = _T_5[_T_5__T_205_addr]; // @[pe.scala 94:49]
  `else
  assign _T_5__T_205_data = _T_5__T_205_addr >= 4'hc ? _RAND_21[127:0] : _T_5[_T_5__T_205_addr]; // @[pe.scala 94:49]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_5__T_78_data = io_to_pes_5_out_bits;
  assign _T_5__T_78_addr = _T_27[3:0];
  assign _T_5__T_78_mask = 1'h1;
  assign _T_5__T_78_en = io_to_pes_5_out_valid;
  assign _T_6__T_207_addr = _T_6__T_207_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_6__T_207_data = _T_6[_T_6__T_207_addr]; // @[pe.scala 94:49]
  `else
  assign _T_6__T_207_data = _T_6__T_207_addr >= 4'hc ? _RAND_25[127:0] : _T_6[_T_6__T_207_addr]; // @[pe.scala 94:49]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_6__T_84_data = io_to_pes_6_out_bits;
  assign _T_6__T_84_addr = _T_28[3:0];
  assign _T_6__T_84_mask = 1'h1;
  assign _T_6__T_84_en = io_to_pes_6_out_valid;
  assign _T_7__T_209_addr = _T_7__T_209_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_7__T_209_data = _T_7[_T_7__T_209_addr]; // @[pe.scala 94:49]
  `else
  assign _T_7__T_209_data = _T_7__T_209_addr >= 4'hc ? _RAND_29[127:0] : _T_7[_T_7__T_209_addr]; // @[pe.scala 94:49]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_7__T_90_data = io_to_pes_7_out_bits;
  assign _T_7__T_90_addr = _T_29[3:0];
  assign _T_7__T_90_mask = 1'h1;
  assign _T_7__T_90_en = io_to_pes_7_out_valid;
  assign _T_8__T_211_addr = _T_8__T_211_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_8__T_211_data = _T_8[_T_8__T_211_addr]; // @[pe.scala 94:49]
  `else
  assign _T_8__T_211_data = _T_8__T_211_addr >= 4'hc ? _RAND_33[127:0] : _T_8[_T_8__T_211_addr]; // @[pe.scala 94:49]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_8__T_96_data = io_to_pes_8_out_bits;
  assign _T_8__T_96_addr = _T_30[3:0];
  assign _T_8__T_96_mask = 1'h1;
  assign _T_8__T_96_en = io_to_pes_8_out_valid;
  assign _T_9__T_213_addr = _T_9__T_213_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_9__T_213_data = _T_9[_T_9__T_213_addr]; // @[pe.scala 94:49]
  `else
  assign _T_9__T_213_data = _T_9__T_213_addr >= 4'hc ? _RAND_37[127:0] : _T_9[_T_9__T_213_addr]; // @[pe.scala 94:49]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_9__T_102_data = io_to_pes_9_out_bits;
  assign _T_9__T_102_addr = _T_31[3:0];
  assign _T_9__T_102_mask = 1'h1;
  assign _T_9__T_102_en = io_to_pes_9_out_valid;
  assign _T_10__T_215_addr = _T_10__T_215_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_10__T_215_data = _T_10[_T_10__T_215_addr]; // @[pe.scala 94:49]
  `else
  assign _T_10__T_215_data = _T_10__T_215_addr >= 4'hc ? _RAND_41[127:0] : _T_10[_T_10__T_215_addr]; // @[pe.scala 94:49]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_10__T_108_data = io_to_pes_10_out_bits;
  assign _T_10__T_108_addr = _T_32[3:0];
  assign _T_10__T_108_mask = 1'h1;
  assign _T_10__T_108_en = io_to_pes_10_out_valid;
  assign _T_11__T_217_addr = _T_11__T_217_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_11__T_217_data = _T_11[_T_11__T_217_addr]; // @[pe.scala 94:49]
  `else
  assign _T_11__T_217_data = _T_11__T_217_addr >= 4'hc ? _RAND_45[127:0] : _T_11[_T_11__T_217_addr]; // @[pe.scala 94:49]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_11__T_114_data = io_to_pes_11_out_bits;
  assign _T_11__T_114_addr = _T_33[3:0];
  assign _T_11__T_114_mask = 1'h1;
  assign _T_11__T_114_en = io_to_pes_11_out_valid;
  assign _T_12__T_219_addr = _T_12__T_219_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_12__T_219_data = _T_12[_T_12__T_219_addr]; // @[pe.scala 94:49]
  `else
  assign _T_12__T_219_data = _T_12__T_219_addr >= 4'hc ? _RAND_49[127:0] : _T_12[_T_12__T_219_addr]; // @[pe.scala 94:49]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_12__T_120_data = io_to_pes_12_out_bits;
  assign _T_12__T_120_addr = _T_34[3:0];
  assign _T_12__T_120_mask = 1'h1;
  assign _T_12__T_120_en = io_to_pes_12_out_valid;
  assign _T_13__T_221_addr = _T_13__T_221_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_13__T_221_data = _T_13[_T_13__T_221_addr]; // @[pe.scala 94:49]
  `else
  assign _T_13__T_221_data = _T_13__T_221_addr >= 4'hc ? _RAND_53[127:0] : _T_13[_T_13__T_221_addr]; // @[pe.scala 94:49]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_13__T_126_data = io_to_pes_13_out_bits;
  assign _T_13__T_126_addr = _T_35[3:0];
  assign _T_13__T_126_mask = 1'h1;
  assign _T_13__T_126_en = io_to_pes_13_out_valid;
  assign _T_14__T_223_addr = _T_14__T_223_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_14__T_223_data = _T_14[_T_14__T_223_addr]; // @[pe.scala 94:49]
  `else
  assign _T_14__T_223_data = _T_14__T_223_addr >= 4'hc ? _RAND_57[127:0] : _T_14[_T_14__T_223_addr]; // @[pe.scala 94:49]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_14__T_132_data = io_to_pes_14_out_bits;
  assign _T_14__T_132_addr = _T_36[3:0];
  assign _T_14__T_132_mask = 1'h1;
  assign _T_14__T_132_en = io_to_pes_14_out_valid;
  assign _T_15__T_225_addr = _T_15__T_225_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_15__T_225_data = _T_15[_T_15__T_225_addr]; // @[pe.scala 94:49]
  `else
  assign _T_15__T_225_data = _T_15__T_225_addr >= 4'hc ? _RAND_61[127:0] : _T_15[_T_15__T_225_addr]; // @[pe.scala 94:49]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_15__T_138_data = io_to_pes_15_out_bits;
  assign _T_15__T_138_addr = _T_37[3:0];
  assign _T_15__T_138_mask = 1'h1;
  assign _T_15__T_138_en = io_to_pes_15_out_valid;
  assign _T_16__T_227_addr = _T_16__T_227_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_16__T_227_data = _T_16[_T_16__T_227_addr]; // @[pe.scala 94:49]
  `else
  assign _T_16__T_227_data = _T_16__T_227_addr >= 4'hc ? _RAND_65[127:0] : _T_16[_T_16__T_227_addr]; // @[pe.scala 94:49]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_16__T_144_data = io_to_pes_16_out_bits;
  assign _T_16__T_144_addr = _T_38[3:0];
  assign _T_16__T_144_mask = 1'h1;
  assign _T_16__T_144_en = io_to_pes_16_out_valid;
  assign _T_17__T_229_addr = _T_17__T_229_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_17__T_229_data = _T_17[_T_17__T_229_addr]; // @[pe.scala 94:49]
  `else
  assign _T_17__T_229_data = _T_17__T_229_addr >= 4'hc ? _RAND_69[127:0] : _T_17[_T_17__T_229_addr]; // @[pe.scala 94:49]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_17__T_150_data = io_to_pes_17_out_bits;
  assign _T_17__T_150_addr = _T_39[3:0];
  assign _T_17__T_150_mask = 1'h1;
  assign _T_17__T_150_en = io_to_pes_17_out_valid;
  assign _T_18__T_231_addr = _T_18__T_231_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_18__T_231_data = _T_18[_T_18__T_231_addr]; // @[pe.scala 94:49]
  `else
  assign _T_18__T_231_data = _T_18__T_231_addr >= 4'hc ? _RAND_73[127:0] : _T_18[_T_18__T_231_addr]; // @[pe.scala 94:49]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_18__T_156_data = io_to_pes_18_out_bits;
  assign _T_18__T_156_addr = _T_40[3:0];
  assign _T_18__T_156_mask = 1'h1;
  assign _T_18__T_156_en = io_to_pes_18_out_valid;
  assign _T_19__T_233_addr = _T_19__T_233_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_19__T_233_data = _T_19[_T_19__T_233_addr]; // @[pe.scala 94:49]
  `else
  assign _T_19__T_233_data = _T_19__T_233_addr >= 4'hc ? _RAND_77[127:0] : _T_19[_T_19__T_233_addr]; // @[pe.scala 94:49]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_19__T_162_data = io_to_pes_19_out_bits;
  assign _T_19__T_162_addr = _T_41[3:0];
  assign _T_19__T_162_mask = 1'h1;
  assign _T_19__T_162_en = io_to_pes_19_out_valid;
  assign _T_20__T_235_addr = _T_20__T_235_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_20__T_235_data = _T_20[_T_20__T_235_addr]; // @[pe.scala 94:49]
  `else
  assign _T_20__T_235_data = _T_20__T_235_addr >= 4'hc ? _RAND_81[127:0] : _T_20[_T_20__T_235_addr]; // @[pe.scala 94:49]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_20__T_168_data = io_to_pes_20_out_bits;
  assign _T_20__T_168_addr = _T_42[3:0];
  assign _T_20__T_168_mask = 1'h1;
  assign _T_20__T_168_en = io_to_pes_20_out_valid;
  assign _T_21__T_237_addr = _T_21__T_237_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_21__T_237_data = _T_21[_T_21__T_237_addr]; // @[pe.scala 94:49]
  `else
  assign _T_21__T_237_data = _T_21__T_237_addr >= 4'hc ? _RAND_85[127:0] : _T_21[_T_21__T_237_addr]; // @[pe.scala 94:49]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_21__T_174_data = io_to_pes_21_out_bits;
  assign _T_21__T_174_addr = _T_43[3:0];
  assign _T_21__T_174_mask = 1'h1;
  assign _T_21__T_174_en = io_to_pes_21_out_valid;
  assign io_to_pes_0_sig_stat2trans = _T_254; // @[pe.scala 142:41]
  assign io_to_pes_1_sig_stat2trans = _T_269; // @[pe.scala 142:41]
  assign io_to_pes_2_sig_stat2trans = _T_284; // @[pe.scala 142:41]
  assign io_to_pes_3_sig_stat2trans = _T_299; // @[pe.scala 142:41]
  assign io_to_pes_4_sig_stat2trans = _T_314; // @[pe.scala 142:41]
  assign io_to_pes_5_sig_stat2trans = _T_329; // @[pe.scala 142:41]
  assign io_to_pes_6_sig_stat2trans = _T_344; // @[pe.scala 142:41]
  assign io_to_pes_7_sig_stat2trans = _T_359; // @[pe.scala 142:41]
  assign io_to_pes_8_sig_stat2trans = _T_374; // @[pe.scala 142:41]
  assign io_to_pes_9_sig_stat2trans = _T_389; // @[pe.scala 142:41]
  assign io_to_pes_10_sig_stat2trans = _T_404; // @[pe.scala 142:41]
  assign io_to_pes_11_sig_stat2trans = _T_419; // @[pe.scala 142:41]
  assign io_to_pes_12_sig_stat2trans = _T_434; // @[pe.scala 142:41]
  assign io_to_pes_13_sig_stat2trans = _T_449; // @[pe.scala 142:41]
  assign io_to_pes_14_sig_stat2trans = _T_464; // @[pe.scala 142:41]
  assign io_to_pes_15_sig_stat2trans = _T_479; // @[pe.scala 142:41]
  assign io_to_pes_16_sig_stat2trans = _T_494; // @[pe.scala 142:41]
  assign io_to_pes_17_sig_stat2trans = _T_509; // @[pe.scala 142:41]
  assign io_to_pes_18_sig_stat2trans = _T_524; // @[pe.scala 142:41]
  assign io_to_pes_19_sig_stat2trans = _T_539; // @[pe.scala 142:41]
  assign io_to_pes_20_sig_stat2trans = _T_554; // @[pe.scala 142:41]
  assign io_to_pes_21_sig_stat2trans = _T_569; // @[pe.scala 142:41]
  assign io_to_mem_valid = _T_44; // @[pe.scala 120:21]
  assign io_to_mem_bits = 5'h15 == _T_46[4:0] ? _T_238_21 : _GEN_157; // @[pe.scala 121:20]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {4{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 12; initvar = initvar+1)
    _T[initvar] = _RAND_0[127:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {4{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T__T_195_en_pipe_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T__T_195_addr_pipe_0 = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_4 = {4{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 12; initvar = initvar+1)
    _T_1[initvar] = _RAND_4[127:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {4{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_1__T_197_en_pipe_0 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_1__T_197_addr_pipe_0 = _RAND_7[3:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_8 = {4{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 12; initvar = initvar+1)
    _T_2[initvar] = _RAND_8[127:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_9 = {4{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_2__T_199_en_pipe_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_2__T_199_addr_pipe_0 = _RAND_11[3:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_12 = {4{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 12; initvar = initvar+1)
    _T_3[initvar] = _RAND_12[127:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_13 = {4{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_3__T_201_en_pipe_0 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_3__T_201_addr_pipe_0 = _RAND_15[3:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_16 = {4{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 12; initvar = initvar+1)
    _T_4[initvar] = _RAND_16[127:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_17 = {4{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_4__T_203_en_pipe_0 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_4__T_203_addr_pipe_0 = _RAND_19[3:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_20 = {4{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 12; initvar = initvar+1)
    _T_5[initvar] = _RAND_20[127:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_21 = {4{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_5__T_205_en_pipe_0 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_5__T_205_addr_pipe_0 = _RAND_23[3:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_24 = {4{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 12; initvar = initvar+1)
    _T_6[initvar] = _RAND_24[127:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_25 = {4{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_6__T_207_en_pipe_0 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_6__T_207_addr_pipe_0 = _RAND_27[3:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_28 = {4{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 12; initvar = initvar+1)
    _T_7[initvar] = _RAND_28[127:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_29 = {4{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_7__T_209_en_pipe_0 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_7__T_209_addr_pipe_0 = _RAND_31[3:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_32 = {4{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 12; initvar = initvar+1)
    _T_8[initvar] = _RAND_32[127:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_33 = {4{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_8__T_211_en_pipe_0 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_8__T_211_addr_pipe_0 = _RAND_35[3:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_36 = {4{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 12; initvar = initvar+1)
    _T_9[initvar] = _RAND_36[127:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_37 = {4{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_9__T_213_en_pipe_0 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_9__T_213_addr_pipe_0 = _RAND_39[3:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_40 = {4{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 12; initvar = initvar+1)
    _T_10[initvar] = _RAND_40[127:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_41 = {4{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_10__T_215_en_pipe_0 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_10__T_215_addr_pipe_0 = _RAND_43[3:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_44 = {4{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 12; initvar = initvar+1)
    _T_11[initvar] = _RAND_44[127:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_45 = {4{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_11__T_217_en_pipe_0 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_11__T_217_addr_pipe_0 = _RAND_47[3:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_48 = {4{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 12; initvar = initvar+1)
    _T_12[initvar] = _RAND_48[127:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_49 = {4{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_12__T_219_en_pipe_0 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_12__T_219_addr_pipe_0 = _RAND_51[3:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_52 = {4{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 12; initvar = initvar+1)
    _T_13[initvar] = _RAND_52[127:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_53 = {4{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T_13__T_221_en_pipe_0 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T_13__T_221_addr_pipe_0 = _RAND_55[3:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_56 = {4{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 12; initvar = initvar+1)
    _T_14[initvar] = _RAND_56[127:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_57 = {4{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T_14__T_223_en_pipe_0 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T_14__T_223_addr_pipe_0 = _RAND_59[3:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_60 = {4{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 12; initvar = initvar+1)
    _T_15[initvar] = _RAND_60[127:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_61 = {4{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T_15__T_225_en_pipe_0 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T_15__T_225_addr_pipe_0 = _RAND_63[3:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_64 = {4{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 12; initvar = initvar+1)
    _T_16[initvar] = _RAND_64[127:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_65 = {4{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _T_16__T_227_en_pipe_0 = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _T_16__T_227_addr_pipe_0 = _RAND_67[3:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_68 = {4{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 12; initvar = initvar+1)
    _T_17[initvar] = _RAND_68[127:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_69 = {4{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _T_17__T_229_en_pipe_0 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _T_17__T_229_addr_pipe_0 = _RAND_71[3:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_72 = {4{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 12; initvar = initvar+1)
    _T_18[initvar] = _RAND_72[127:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_73 = {4{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _T_18__T_231_en_pipe_0 = _RAND_74[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _T_18__T_231_addr_pipe_0 = _RAND_75[3:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_76 = {4{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 12; initvar = initvar+1)
    _T_19[initvar] = _RAND_76[127:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_77 = {4{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  _T_19__T_233_en_pipe_0 = _RAND_78[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  _T_19__T_233_addr_pipe_0 = _RAND_79[3:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_80 = {4{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 12; initvar = initvar+1)
    _T_20[initvar] = _RAND_80[127:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_81 = {4{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _T_20__T_235_en_pipe_0 = _RAND_82[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _T_20__T_235_addr_pipe_0 = _RAND_83[3:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_84 = {4{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 12; initvar = initvar+1)
    _T_21[initvar] = _RAND_84[127:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_85 = {4{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _T_21__T_237_en_pipe_0 = _RAND_86[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  _T_21__T_237_addr_pipe_0 = _RAND_87[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  _T_22 = _RAND_88[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  _T_23 = _RAND_89[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  _T_24 = _RAND_90[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  _T_25 = _RAND_91[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  _T_26 = _RAND_92[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  _T_27 = _RAND_93[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _T_28 = _RAND_94[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  _T_29 = _RAND_95[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  _T_30 = _RAND_96[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  _T_31 = _RAND_97[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  _T_32 = _RAND_98[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  _T_33 = _RAND_99[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  _T_34 = _RAND_100[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  _T_35 = _RAND_101[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  _T_36 = _RAND_102[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  _T_37 = _RAND_103[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  _T_38 = _RAND_104[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  _T_39 = _RAND_105[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  _T_40 = _RAND_106[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  _T_41 = _RAND_107[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  _T_42 = _RAND_108[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  _T_43 = _RAND_109[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  _T_44 = _RAND_110[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  _T_45 = _RAND_111[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  _T_46 = _RAND_112[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  _T_240 = _RAND_113[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  _T_241 = _RAND_114[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  _T_242 = _RAND_115[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  _T_243 = _RAND_116[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  _T_244 = _RAND_117[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  _T_245 = _RAND_118[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  _T_246 = _RAND_119[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  _T_247 = _RAND_120[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  _T_248 = _RAND_121[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  _T_249 = _RAND_122[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  _T_250 = _RAND_123[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  _T_251 = _RAND_124[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  _T_252 = _RAND_125[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  _T_253 = _RAND_126[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  _T_254 = _RAND_127[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  _T_255 = _RAND_128[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  _T_256 = _RAND_129[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  _T_257 = _RAND_130[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  _T_258 = _RAND_131[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  _T_259 = _RAND_132[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  _T_260 = _RAND_133[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  _T_261 = _RAND_134[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  _T_262 = _RAND_135[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  _T_263 = _RAND_136[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  _T_264 = _RAND_137[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  _T_265 = _RAND_138[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  _T_266 = _RAND_139[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  _T_267 = _RAND_140[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  _T_268 = _RAND_141[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  _T_269 = _RAND_142[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  _T_270 = _RAND_143[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  _T_271 = _RAND_144[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  _T_272 = _RAND_145[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  _T_273 = _RAND_146[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  _T_274 = _RAND_147[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  _T_275 = _RAND_148[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  _T_276 = _RAND_149[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  _T_277 = _RAND_150[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  _T_278 = _RAND_151[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  _T_279 = _RAND_152[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  _T_280 = _RAND_153[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  _T_281 = _RAND_154[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  _T_282 = _RAND_155[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  _T_283 = _RAND_156[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  _T_284 = _RAND_157[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  _T_285 = _RAND_158[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  _T_286 = _RAND_159[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  _T_287 = _RAND_160[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  _T_288 = _RAND_161[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  _T_289 = _RAND_162[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  _T_290 = _RAND_163[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  _T_291 = _RAND_164[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  _T_292 = _RAND_165[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  _T_293 = _RAND_166[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  _T_294 = _RAND_167[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  _T_295 = _RAND_168[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  _T_296 = _RAND_169[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  _T_297 = _RAND_170[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  _T_298 = _RAND_171[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  _T_299 = _RAND_172[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  _T_300 = _RAND_173[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  _T_301 = _RAND_174[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  _T_302 = _RAND_175[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  _T_303 = _RAND_176[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  _T_304 = _RAND_177[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  _T_305 = _RAND_178[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  _T_306 = _RAND_179[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  _T_307 = _RAND_180[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  _T_308 = _RAND_181[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  _T_309 = _RAND_182[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  _T_310 = _RAND_183[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  _T_311 = _RAND_184[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  _T_312 = _RAND_185[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  _T_313 = _RAND_186[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  _T_314 = _RAND_187[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  _T_315 = _RAND_188[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  _T_316 = _RAND_189[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  _T_317 = _RAND_190[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  _T_318 = _RAND_191[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  _T_319 = _RAND_192[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  _T_320 = _RAND_193[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  _T_321 = _RAND_194[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  _T_322 = _RAND_195[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  _T_323 = _RAND_196[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  _T_324 = _RAND_197[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  _T_325 = _RAND_198[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  _T_326 = _RAND_199[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  _T_327 = _RAND_200[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  _T_328 = _RAND_201[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  _T_329 = _RAND_202[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  _T_330 = _RAND_203[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  _T_331 = _RAND_204[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  _T_332 = _RAND_205[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  _T_333 = _RAND_206[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  _T_334 = _RAND_207[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  _T_335 = _RAND_208[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  _T_336 = _RAND_209[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  _T_337 = _RAND_210[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  _T_338 = _RAND_211[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{`RANDOM}};
  _T_339 = _RAND_212[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{`RANDOM}};
  _T_340 = _RAND_213[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{`RANDOM}};
  _T_341 = _RAND_214[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{`RANDOM}};
  _T_342 = _RAND_215[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{`RANDOM}};
  _T_343 = _RAND_216[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{`RANDOM}};
  _T_344 = _RAND_217[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{`RANDOM}};
  _T_345 = _RAND_218[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{`RANDOM}};
  _T_346 = _RAND_219[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{`RANDOM}};
  _T_347 = _RAND_220[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{`RANDOM}};
  _T_348 = _RAND_221[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{`RANDOM}};
  _T_349 = _RAND_222[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{`RANDOM}};
  _T_350 = _RAND_223[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{`RANDOM}};
  _T_351 = _RAND_224[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{`RANDOM}};
  _T_352 = _RAND_225[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{`RANDOM}};
  _T_353 = _RAND_226[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{`RANDOM}};
  _T_354 = _RAND_227[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{`RANDOM}};
  _T_355 = _RAND_228[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{`RANDOM}};
  _T_356 = _RAND_229[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{`RANDOM}};
  _T_357 = _RAND_230[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{`RANDOM}};
  _T_358 = _RAND_231[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{`RANDOM}};
  _T_359 = _RAND_232[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{`RANDOM}};
  _T_360 = _RAND_233[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{`RANDOM}};
  _T_361 = _RAND_234[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{`RANDOM}};
  _T_362 = _RAND_235[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{`RANDOM}};
  _T_363 = _RAND_236[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{`RANDOM}};
  _T_364 = _RAND_237[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{`RANDOM}};
  _T_365 = _RAND_238[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{`RANDOM}};
  _T_366 = _RAND_239[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{`RANDOM}};
  _T_367 = _RAND_240[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{`RANDOM}};
  _T_368 = _RAND_241[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{`RANDOM}};
  _T_369 = _RAND_242[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{`RANDOM}};
  _T_370 = _RAND_243[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{`RANDOM}};
  _T_371 = _RAND_244[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{`RANDOM}};
  _T_372 = _RAND_245[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{`RANDOM}};
  _T_373 = _RAND_246[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{`RANDOM}};
  _T_374 = _RAND_247[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{`RANDOM}};
  _T_375 = _RAND_248[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{`RANDOM}};
  _T_376 = _RAND_249[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{`RANDOM}};
  _T_377 = _RAND_250[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{`RANDOM}};
  _T_378 = _RAND_251[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{`RANDOM}};
  _T_379 = _RAND_252[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{`RANDOM}};
  _T_380 = _RAND_253[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{`RANDOM}};
  _T_381 = _RAND_254[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{`RANDOM}};
  _T_382 = _RAND_255[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{`RANDOM}};
  _T_383 = _RAND_256[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{`RANDOM}};
  _T_384 = _RAND_257[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_258 = {1{`RANDOM}};
  _T_385 = _RAND_258[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_259 = {1{`RANDOM}};
  _T_386 = _RAND_259[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_260 = {1{`RANDOM}};
  _T_387 = _RAND_260[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_261 = {1{`RANDOM}};
  _T_388 = _RAND_261[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_262 = {1{`RANDOM}};
  _T_389 = _RAND_262[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_263 = {1{`RANDOM}};
  _T_390 = _RAND_263[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_264 = {1{`RANDOM}};
  _T_391 = _RAND_264[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_265 = {1{`RANDOM}};
  _T_392 = _RAND_265[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_266 = {1{`RANDOM}};
  _T_393 = _RAND_266[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_267 = {1{`RANDOM}};
  _T_394 = _RAND_267[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_268 = {1{`RANDOM}};
  _T_395 = _RAND_268[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_269 = {1{`RANDOM}};
  _T_396 = _RAND_269[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_270 = {1{`RANDOM}};
  _T_397 = _RAND_270[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_271 = {1{`RANDOM}};
  _T_398 = _RAND_271[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_272 = {1{`RANDOM}};
  _T_399 = _RAND_272[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_273 = {1{`RANDOM}};
  _T_400 = _RAND_273[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_274 = {1{`RANDOM}};
  _T_401 = _RAND_274[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_275 = {1{`RANDOM}};
  _T_402 = _RAND_275[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_276 = {1{`RANDOM}};
  _T_403 = _RAND_276[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_277 = {1{`RANDOM}};
  _T_404 = _RAND_277[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_278 = {1{`RANDOM}};
  _T_405 = _RAND_278[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_279 = {1{`RANDOM}};
  _T_406 = _RAND_279[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_280 = {1{`RANDOM}};
  _T_407 = _RAND_280[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_281 = {1{`RANDOM}};
  _T_408 = _RAND_281[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_282 = {1{`RANDOM}};
  _T_409 = _RAND_282[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_283 = {1{`RANDOM}};
  _T_410 = _RAND_283[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_284 = {1{`RANDOM}};
  _T_411 = _RAND_284[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_285 = {1{`RANDOM}};
  _T_412 = _RAND_285[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_286 = {1{`RANDOM}};
  _T_413 = _RAND_286[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_287 = {1{`RANDOM}};
  _T_414 = _RAND_287[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_288 = {1{`RANDOM}};
  _T_415 = _RAND_288[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_289 = {1{`RANDOM}};
  _T_416 = _RAND_289[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_290 = {1{`RANDOM}};
  _T_417 = _RAND_290[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_291 = {1{`RANDOM}};
  _T_418 = _RAND_291[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_292 = {1{`RANDOM}};
  _T_419 = _RAND_292[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_293 = {1{`RANDOM}};
  _T_420 = _RAND_293[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_294 = {1{`RANDOM}};
  _T_421 = _RAND_294[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_295 = {1{`RANDOM}};
  _T_422 = _RAND_295[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_296 = {1{`RANDOM}};
  _T_423 = _RAND_296[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_297 = {1{`RANDOM}};
  _T_424 = _RAND_297[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_298 = {1{`RANDOM}};
  _T_425 = _RAND_298[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_299 = {1{`RANDOM}};
  _T_426 = _RAND_299[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_300 = {1{`RANDOM}};
  _T_427 = _RAND_300[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_301 = {1{`RANDOM}};
  _T_428 = _RAND_301[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_302 = {1{`RANDOM}};
  _T_429 = _RAND_302[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_303 = {1{`RANDOM}};
  _T_430 = _RAND_303[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_304 = {1{`RANDOM}};
  _T_431 = _RAND_304[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_305 = {1{`RANDOM}};
  _T_432 = _RAND_305[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_306 = {1{`RANDOM}};
  _T_433 = _RAND_306[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_307 = {1{`RANDOM}};
  _T_434 = _RAND_307[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_308 = {1{`RANDOM}};
  _T_435 = _RAND_308[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_309 = {1{`RANDOM}};
  _T_436 = _RAND_309[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_310 = {1{`RANDOM}};
  _T_437 = _RAND_310[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_311 = {1{`RANDOM}};
  _T_438 = _RAND_311[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_312 = {1{`RANDOM}};
  _T_439 = _RAND_312[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_313 = {1{`RANDOM}};
  _T_440 = _RAND_313[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_314 = {1{`RANDOM}};
  _T_441 = _RAND_314[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_315 = {1{`RANDOM}};
  _T_442 = _RAND_315[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_316 = {1{`RANDOM}};
  _T_443 = _RAND_316[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_317 = {1{`RANDOM}};
  _T_444 = _RAND_317[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_318 = {1{`RANDOM}};
  _T_445 = _RAND_318[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_319 = {1{`RANDOM}};
  _T_446 = _RAND_319[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_320 = {1{`RANDOM}};
  _T_447 = _RAND_320[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_321 = {1{`RANDOM}};
  _T_448 = _RAND_321[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_322 = {1{`RANDOM}};
  _T_449 = _RAND_322[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_323 = {1{`RANDOM}};
  _T_450 = _RAND_323[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_324 = {1{`RANDOM}};
  _T_451 = _RAND_324[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_325 = {1{`RANDOM}};
  _T_452 = _RAND_325[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_326 = {1{`RANDOM}};
  _T_453 = _RAND_326[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_327 = {1{`RANDOM}};
  _T_454 = _RAND_327[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_328 = {1{`RANDOM}};
  _T_455 = _RAND_328[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_329 = {1{`RANDOM}};
  _T_456 = _RAND_329[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_330 = {1{`RANDOM}};
  _T_457 = _RAND_330[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_331 = {1{`RANDOM}};
  _T_458 = _RAND_331[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_332 = {1{`RANDOM}};
  _T_459 = _RAND_332[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_333 = {1{`RANDOM}};
  _T_460 = _RAND_333[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_334 = {1{`RANDOM}};
  _T_461 = _RAND_334[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_335 = {1{`RANDOM}};
  _T_462 = _RAND_335[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_336 = {1{`RANDOM}};
  _T_463 = _RAND_336[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_337 = {1{`RANDOM}};
  _T_464 = _RAND_337[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_338 = {1{`RANDOM}};
  _T_465 = _RAND_338[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_339 = {1{`RANDOM}};
  _T_466 = _RAND_339[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_340 = {1{`RANDOM}};
  _T_467 = _RAND_340[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_341 = {1{`RANDOM}};
  _T_468 = _RAND_341[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_342 = {1{`RANDOM}};
  _T_469 = _RAND_342[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_343 = {1{`RANDOM}};
  _T_470 = _RAND_343[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_344 = {1{`RANDOM}};
  _T_471 = _RAND_344[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_345 = {1{`RANDOM}};
  _T_472 = _RAND_345[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_346 = {1{`RANDOM}};
  _T_473 = _RAND_346[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_347 = {1{`RANDOM}};
  _T_474 = _RAND_347[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_348 = {1{`RANDOM}};
  _T_475 = _RAND_348[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_349 = {1{`RANDOM}};
  _T_476 = _RAND_349[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_350 = {1{`RANDOM}};
  _T_477 = _RAND_350[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_351 = {1{`RANDOM}};
  _T_478 = _RAND_351[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_352 = {1{`RANDOM}};
  _T_479 = _RAND_352[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_353 = {1{`RANDOM}};
  _T_480 = _RAND_353[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_354 = {1{`RANDOM}};
  _T_481 = _RAND_354[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_355 = {1{`RANDOM}};
  _T_482 = _RAND_355[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_356 = {1{`RANDOM}};
  _T_483 = _RAND_356[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_357 = {1{`RANDOM}};
  _T_484 = _RAND_357[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_358 = {1{`RANDOM}};
  _T_485 = _RAND_358[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_359 = {1{`RANDOM}};
  _T_486 = _RAND_359[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_360 = {1{`RANDOM}};
  _T_487 = _RAND_360[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_361 = {1{`RANDOM}};
  _T_488 = _RAND_361[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_362 = {1{`RANDOM}};
  _T_489 = _RAND_362[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_363 = {1{`RANDOM}};
  _T_490 = _RAND_363[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_364 = {1{`RANDOM}};
  _T_491 = _RAND_364[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_365 = {1{`RANDOM}};
  _T_492 = _RAND_365[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_366 = {1{`RANDOM}};
  _T_493 = _RAND_366[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_367 = {1{`RANDOM}};
  _T_494 = _RAND_367[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_368 = {1{`RANDOM}};
  _T_495 = _RAND_368[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_369 = {1{`RANDOM}};
  _T_496 = _RAND_369[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_370 = {1{`RANDOM}};
  _T_497 = _RAND_370[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_371 = {1{`RANDOM}};
  _T_498 = _RAND_371[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_372 = {1{`RANDOM}};
  _T_499 = _RAND_372[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_373 = {1{`RANDOM}};
  _T_500 = _RAND_373[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_374 = {1{`RANDOM}};
  _T_501 = _RAND_374[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_375 = {1{`RANDOM}};
  _T_502 = _RAND_375[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_376 = {1{`RANDOM}};
  _T_503 = _RAND_376[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_377 = {1{`RANDOM}};
  _T_504 = _RAND_377[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_378 = {1{`RANDOM}};
  _T_505 = _RAND_378[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_379 = {1{`RANDOM}};
  _T_506 = _RAND_379[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_380 = {1{`RANDOM}};
  _T_507 = _RAND_380[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_381 = {1{`RANDOM}};
  _T_508 = _RAND_381[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_382 = {1{`RANDOM}};
  _T_509 = _RAND_382[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_383 = {1{`RANDOM}};
  _T_510 = _RAND_383[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_384 = {1{`RANDOM}};
  _T_511 = _RAND_384[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_385 = {1{`RANDOM}};
  _T_512 = _RAND_385[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_386 = {1{`RANDOM}};
  _T_513 = _RAND_386[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_387 = {1{`RANDOM}};
  _T_514 = _RAND_387[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_388 = {1{`RANDOM}};
  _T_515 = _RAND_388[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_389 = {1{`RANDOM}};
  _T_516 = _RAND_389[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_390 = {1{`RANDOM}};
  _T_517 = _RAND_390[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_391 = {1{`RANDOM}};
  _T_518 = _RAND_391[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_392 = {1{`RANDOM}};
  _T_519 = _RAND_392[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_393 = {1{`RANDOM}};
  _T_520 = _RAND_393[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_394 = {1{`RANDOM}};
  _T_521 = _RAND_394[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_395 = {1{`RANDOM}};
  _T_522 = _RAND_395[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_396 = {1{`RANDOM}};
  _T_523 = _RAND_396[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_397 = {1{`RANDOM}};
  _T_524 = _RAND_397[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_398 = {1{`RANDOM}};
  _T_525 = _RAND_398[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_399 = {1{`RANDOM}};
  _T_526 = _RAND_399[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_400 = {1{`RANDOM}};
  _T_527 = _RAND_400[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_401 = {1{`RANDOM}};
  _T_528 = _RAND_401[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_402 = {1{`RANDOM}};
  _T_529 = _RAND_402[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_403 = {1{`RANDOM}};
  _T_530 = _RAND_403[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_404 = {1{`RANDOM}};
  _T_531 = _RAND_404[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_405 = {1{`RANDOM}};
  _T_532 = _RAND_405[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_406 = {1{`RANDOM}};
  _T_533 = _RAND_406[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_407 = {1{`RANDOM}};
  _T_534 = _RAND_407[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_408 = {1{`RANDOM}};
  _T_535 = _RAND_408[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_409 = {1{`RANDOM}};
  _T_536 = _RAND_409[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_410 = {1{`RANDOM}};
  _T_537 = _RAND_410[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_411 = {1{`RANDOM}};
  _T_538 = _RAND_411[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_412 = {1{`RANDOM}};
  _T_539 = _RAND_412[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_413 = {1{`RANDOM}};
  _T_540 = _RAND_413[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_414 = {1{`RANDOM}};
  _T_541 = _RAND_414[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_415 = {1{`RANDOM}};
  _T_542 = _RAND_415[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_416 = {1{`RANDOM}};
  _T_543 = _RAND_416[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_417 = {1{`RANDOM}};
  _T_544 = _RAND_417[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_418 = {1{`RANDOM}};
  _T_545 = _RAND_418[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_419 = {1{`RANDOM}};
  _T_546 = _RAND_419[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_420 = {1{`RANDOM}};
  _T_547 = _RAND_420[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_421 = {1{`RANDOM}};
  _T_548 = _RAND_421[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_422 = {1{`RANDOM}};
  _T_549 = _RAND_422[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_423 = {1{`RANDOM}};
  _T_550 = _RAND_423[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_424 = {1{`RANDOM}};
  _T_551 = _RAND_424[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_425 = {1{`RANDOM}};
  _T_552 = _RAND_425[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_426 = {1{`RANDOM}};
  _T_553 = _RAND_426[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_427 = {1{`RANDOM}};
  _T_554 = _RAND_427[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_428 = {1{`RANDOM}};
  _T_555 = _RAND_428[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_429 = {1{`RANDOM}};
  _T_556 = _RAND_429[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_430 = {1{`RANDOM}};
  _T_557 = _RAND_430[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_431 = {1{`RANDOM}};
  _T_558 = _RAND_431[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_432 = {1{`RANDOM}};
  _T_559 = _RAND_432[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_433 = {1{`RANDOM}};
  _T_560 = _RAND_433[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_434 = {1{`RANDOM}};
  _T_561 = _RAND_434[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_435 = {1{`RANDOM}};
  _T_562 = _RAND_435[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_436 = {1{`RANDOM}};
  _T_563 = _RAND_436[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_437 = {1{`RANDOM}};
  _T_564 = _RAND_437[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_438 = {1{`RANDOM}};
  _T_565 = _RAND_438[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_439 = {1{`RANDOM}};
  _T_566 = _RAND_439[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_440 = {1{`RANDOM}};
  _T_567 = _RAND_440[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_441 = {1{`RANDOM}};
  _T_568 = _RAND_441[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_442 = {1{`RANDOM}};
  _T_569 = _RAND_442[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T__T_48_en & _T__T_48_mask) begin
      _T[_T__T_48_addr] <= _T__T_48_data; // @[pe.scala 94:49]
    end
    _T__T_195_en_pipe_0 <= 1'h1;
    _T__T_195_addr_pipe_0 <= _T_45[3:0];
    if(_T_1__T_54_en & _T_1__T_54_mask) begin
      _T_1[_T_1__T_54_addr] <= _T_1__T_54_data; // @[pe.scala 94:49]
    end
    _T_1__T_197_en_pipe_0 <= 1'h1;
    _T_1__T_197_addr_pipe_0 <= _T_45[3:0];
    if(_T_2__T_60_en & _T_2__T_60_mask) begin
      _T_2[_T_2__T_60_addr] <= _T_2__T_60_data; // @[pe.scala 94:49]
    end
    _T_2__T_199_en_pipe_0 <= 1'h1;
    _T_2__T_199_addr_pipe_0 <= _T_45[3:0];
    if(_T_3__T_66_en & _T_3__T_66_mask) begin
      _T_3[_T_3__T_66_addr] <= _T_3__T_66_data; // @[pe.scala 94:49]
    end
    _T_3__T_201_en_pipe_0 <= 1'h1;
    _T_3__T_201_addr_pipe_0 <= _T_45[3:0];
    if(_T_4__T_72_en & _T_4__T_72_mask) begin
      _T_4[_T_4__T_72_addr] <= _T_4__T_72_data; // @[pe.scala 94:49]
    end
    _T_4__T_203_en_pipe_0 <= 1'h1;
    _T_4__T_203_addr_pipe_0 <= _T_45[3:0];
    if(_T_5__T_78_en & _T_5__T_78_mask) begin
      _T_5[_T_5__T_78_addr] <= _T_5__T_78_data; // @[pe.scala 94:49]
    end
    _T_5__T_205_en_pipe_0 <= 1'h1;
    _T_5__T_205_addr_pipe_0 <= _T_45[3:0];
    if(_T_6__T_84_en & _T_6__T_84_mask) begin
      _T_6[_T_6__T_84_addr] <= _T_6__T_84_data; // @[pe.scala 94:49]
    end
    _T_6__T_207_en_pipe_0 <= 1'h1;
    _T_6__T_207_addr_pipe_0 <= _T_45[3:0];
    if(_T_7__T_90_en & _T_7__T_90_mask) begin
      _T_7[_T_7__T_90_addr] <= _T_7__T_90_data; // @[pe.scala 94:49]
    end
    _T_7__T_209_en_pipe_0 <= 1'h1;
    _T_7__T_209_addr_pipe_0 <= _T_45[3:0];
    if(_T_8__T_96_en & _T_8__T_96_mask) begin
      _T_8[_T_8__T_96_addr] <= _T_8__T_96_data; // @[pe.scala 94:49]
    end
    _T_8__T_211_en_pipe_0 <= 1'h1;
    _T_8__T_211_addr_pipe_0 <= _T_45[3:0];
    if(_T_9__T_102_en & _T_9__T_102_mask) begin
      _T_9[_T_9__T_102_addr] <= _T_9__T_102_data; // @[pe.scala 94:49]
    end
    _T_9__T_213_en_pipe_0 <= 1'h1;
    _T_9__T_213_addr_pipe_0 <= _T_45[3:0];
    if(_T_10__T_108_en & _T_10__T_108_mask) begin
      _T_10[_T_10__T_108_addr] <= _T_10__T_108_data; // @[pe.scala 94:49]
    end
    _T_10__T_215_en_pipe_0 <= 1'h1;
    _T_10__T_215_addr_pipe_0 <= _T_45[3:0];
    if(_T_11__T_114_en & _T_11__T_114_mask) begin
      _T_11[_T_11__T_114_addr] <= _T_11__T_114_data; // @[pe.scala 94:49]
    end
    _T_11__T_217_en_pipe_0 <= 1'h1;
    _T_11__T_217_addr_pipe_0 <= _T_45[3:0];
    if(_T_12__T_120_en & _T_12__T_120_mask) begin
      _T_12[_T_12__T_120_addr] <= _T_12__T_120_data; // @[pe.scala 94:49]
    end
    _T_12__T_219_en_pipe_0 <= 1'h1;
    _T_12__T_219_addr_pipe_0 <= _T_45[3:0];
    if(_T_13__T_126_en & _T_13__T_126_mask) begin
      _T_13[_T_13__T_126_addr] <= _T_13__T_126_data; // @[pe.scala 94:49]
    end
    _T_13__T_221_en_pipe_0 <= 1'h1;
    _T_13__T_221_addr_pipe_0 <= _T_45[3:0];
    if(_T_14__T_132_en & _T_14__T_132_mask) begin
      _T_14[_T_14__T_132_addr] <= _T_14__T_132_data; // @[pe.scala 94:49]
    end
    _T_14__T_223_en_pipe_0 <= 1'h1;
    _T_14__T_223_addr_pipe_0 <= _T_45[3:0];
    if(_T_15__T_138_en & _T_15__T_138_mask) begin
      _T_15[_T_15__T_138_addr] <= _T_15__T_138_data; // @[pe.scala 94:49]
    end
    _T_15__T_225_en_pipe_0 <= 1'h1;
    _T_15__T_225_addr_pipe_0 <= _T_45[3:0];
    if(_T_16__T_144_en & _T_16__T_144_mask) begin
      _T_16[_T_16__T_144_addr] <= _T_16__T_144_data; // @[pe.scala 94:49]
    end
    _T_16__T_227_en_pipe_0 <= 1'h1;
    _T_16__T_227_addr_pipe_0 <= _T_45[3:0];
    if(_T_17__T_150_en & _T_17__T_150_mask) begin
      _T_17[_T_17__T_150_addr] <= _T_17__T_150_data; // @[pe.scala 94:49]
    end
    _T_17__T_229_en_pipe_0 <= 1'h1;
    _T_17__T_229_addr_pipe_0 <= _T_45[3:0];
    if(_T_18__T_156_en & _T_18__T_156_mask) begin
      _T_18[_T_18__T_156_addr] <= _T_18__T_156_data; // @[pe.scala 94:49]
    end
    _T_18__T_231_en_pipe_0 <= 1'h1;
    _T_18__T_231_addr_pipe_0 <= _T_45[3:0];
    if(_T_19__T_162_en & _T_19__T_162_mask) begin
      _T_19[_T_19__T_162_addr] <= _T_19__T_162_data; // @[pe.scala 94:49]
    end
    _T_19__T_233_en_pipe_0 <= 1'h1;
    _T_19__T_233_addr_pipe_0 <= _T_45[3:0];
    if(_T_20__T_168_en & _T_20__T_168_mask) begin
      _T_20[_T_20__T_168_addr] <= _T_20__T_168_data; // @[pe.scala 94:49]
    end
    _T_20__T_235_en_pipe_0 <= 1'h1;
    _T_20__T_235_addr_pipe_0 <= _T_45[3:0];
    if(_T_21__T_174_en & _T_21__T_174_mask) begin
      _T_21[_T_21__T_174_addr] <= _T_21__T_174_data; // @[pe.scala 94:49]
    end
    _T_21__T_237_en_pipe_0 <= 1'h1;
    _T_21__T_237_addr_pipe_0 <= _T_45[3:0];
    if (reset) begin
      _T_22 <= 5'h0;
    end else if (io_to_pes_0_out_valid) begin
      if (_T_49) begin
        _T_22 <= 5'h0;
      end else begin
        _T_22 <= _T_51;
      end
    end
    if (reset) begin
      _T_23 <= 5'h0;
    end else if (io_to_pes_1_out_valid) begin
      if (_T_55) begin
        _T_23 <= 5'h0;
      end else begin
        _T_23 <= _T_57;
      end
    end
    if (reset) begin
      _T_24 <= 5'h0;
    end else if (io_to_pes_2_out_valid) begin
      if (_T_61) begin
        _T_24 <= 5'h0;
      end else begin
        _T_24 <= _T_63;
      end
    end
    if (reset) begin
      _T_25 <= 5'h0;
    end else if (io_to_pes_3_out_valid) begin
      if (_T_67) begin
        _T_25 <= 5'h0;
      end else begin
        _T_25 <= _T_69;
      end
    end
    if (reset) begin
      _T_26 <= 5'h0;
    end else if (io_to_pes_4_out_valid) begin
      if (_T_73) begin
        _T_26 <= 5'h0;
      end else begin
        _T_26 <= _T_75;
      end
    end
    if (reset) begin
      _T_27 <= 5'h0;
    end else if (io_to_pes_5_out_valid) begin
      if (_T_79) begin
        _T_27 <= 5'h0;
      end else begin
        _T_27 <= _T_81;
      end
    end
    if (reset) begin
      _T_28 <= 5'h0;
    end else if (io_to_pes_6_out_valid) begin
      if (_T_85) begin
        _T_28 <= 5'h0;
      end else begin
        _T_28 <= _T_87;
      end
    end
    if (reset) begin
      _T_29 <= 5'h0;
    end else if (io_to_pes_7_out_valid) begin
      if (_T_91) begin
        _T_29 <= 5'h0;
      end else begin
        _T_29 <= _T_93;
      end
    end
    if (reset) begin
      _T_30 <= 5'h0;
    end else if (io_to_pes_8_out_valid) begin
      if (_T_97) begin
        _T_30 <= 5'h0;
      end else begin
        _T_30 <= _T_99;
      end
    end
    if (reset) begin
      _T_31 <= 5'h0;
    end else if (io_to_pes_9_out_valid) begin
      if (_T_103) begin
        _T_31 <= 5'h0;
      end else begin
        _T_31 <= _T_105;
      end
    end
    if (reset) begin
      _T_32 <= 5'h0;
    end else if (io_to_pes_10_out_valid) begin
      if (_T_109) begin
        _T_32 <= 5'h0;
      end else begin
        _T_32 <= _T_111;
      end
    end
    if (reset) begin
      _T_33 <= 5'h0;
    end else if (io_to_pes_11_out_valid) begin
      if (_T_115) begin
        _T_33 <= 5'h0;
      end else begin
        _T_33 <= _T_117;
      end
    end
    if (reset) begin
      _T_34 <= 5'h0;
    end else if (io_to_pes_12_out_valid) begin
      if (_T_121) begin
        _T_34 <= 5'h0;
      end else begin
        _T_34 <= _T_123;
      end
    end
    if (reset) begin
      _T_35 <= 5'h0;
    end else if (io_to_pes_13_out_valid) begin
      if (_T_127) begin
        _T_35 <= 5'h0;
      end else begin
        _T_35 <= _T_129;
      end
    end
    if (reset) begin
      _T_36 <= 5'h0;
    end else if (io_to_pes_14_out_valid) begin
      if (_T_133) begin
        _T_36 <= 5'h0;
      end else begin
        _T_36 <= _T_135;
      end
    end
    if (reset) begin
      _T_37 <= 5'h0;
    end else if (io_to_pes_15_out_valid) begin
      if (_T_139) begin
        _T_37 <= 5'h0;
      end else begin
        _T_37 <= _T_141;
      end
    end
    if (reset) begin
      _T_38 <= 5'h0;
    end else if (io_to_pes_16_out_valid) begin
      if (_T_145) begin
        _T_38 <= 5'h0;
      end else begin
        _T_38 <= _T_147;
      end
    end
    if (reset) begin
      _T_39 <= 5'h0;
    end else if (io_to_pes_17_out_valid) begin
      if (_T_151) begin
        _T_39 <= 5'h0;
      end else begin
        _T_39 <= _T_153;
      end
    end
    if (reset) begin
      _T_40 <= 5'h0;
    end else if (io_to_pes_18_out_valid) begin
      if (_T_157) begin
        _T_40 <= 5'h0;
      end else begin
        _T_40 <= _T_159;
      end
    end
    if (reset) begin
      _T_41 <= 5'h0;
    end else if (io_to_pes_19_out_valid) begin
      if (_T_163) begin
        _T_41 <= 5'h0;
      end else begin
        _T_41 <= _T_165;
      end
    end
    if (reset) begin
      _T_42 <= 5'h0;
    end else if (io_to_pes_20_out_valid) begin
      if (_T_169) begin
        _T_42 <= 5'h0;
      end else begin
        _T_42 <= _T_171;
      end
    end
    if (reset) begin
      _T_43 <= 5'h0;
    end else if (io_to_pes_21_out_valid) begin
      if (_T_175) begin
        _T_43 <= 5'h0;
      end else begin
        _T_43 <= _T_177;
      end
    end
    if (reset) begin
      _T_44 <= 1'h0;
    end else if (_T_44) begin
      if (_T_193) begin
        _T_44 <= 1'h0;
      end else begin
        _T_44 <= _GEN_132;
      end
    end else begin
      _T_44 <= _GEN_132;
    end
    if (reset) begin
      _T_45 <= 10'h0;
    end else if (_T_44) begin
      if (_T_181) begin
        _T_45 <= 10'h0;
      end else begin
        _T_45 <= _T_183;
      end
    end
    if (reset) begin
      _T_46 <= 10'h0;
    end else if (_T_44) begin
      if (_T_181) begin
        if (_T_186) begin
          _T_46 <= 10'h0;
        end else begin
          _T_46 <= _T_188;
        end
      end
    end
    _T_240 <= io_sig_stat2trans;
    _T_241 <= _T_240;
    _T_242 <= _T_241;
    _T_243 <= _T_242;
    _T_244 <= _T_243;
    _T_245 <= _T_244;
    _T_246 <= _T_245;
    _T_247 <= _T_246;
    _T_248 <= _T_247;
    _T_249 <= _T_248;
    _T_250 <= _T_249;
    _T_251 <= _T_250;
    _T_252 <= _T_251;
    _T_253 <= _T_252;
    _T_254 <= _T_253;
    _T_255 <= io_sig_stat2trans;
    _T_256 <= _T_255;
    _T_257 <= _T_256;
    _T_258 <= _T_257;
    _T_259 <= _T_258;
    _T_260 <= _T_259;
    _T_261 <= _T_260;
    _T_262 <= _T_261;
    _T_263 <= _T_262;
    _T_264 <= _T_263;
    _T_265 <= _T_264;
    _T_266 <= _T_265;
    _T_267 <= _T_266;
    _T_268 <= _T_267;
    _T_269 <= _T_268;
    _T_270 <= io_sig_stat2trans;
    _T_271 <= _T_270;
    _T_272 <= _T_271;
    _T_273 <= _T_272;
    _T_274 <= _T_273;
    _T_275 <= _T_274;
    _T_276 <= _T_275;
    _T_277 <= _T_276;
    _T_278 <= _T_277;
    _T_279 <= _T_278;
    _T_280 <= _T_279;
    _T_281 <= _T_280;
    _T_282 <= _T_281;
    _T_283 <= _T_282;
    _T_284 <= _T_283;
    _T_285 <= io_sig_stat2trans;
    _T_286 <= _T_285;
    _T_287 <= _T_286;
    _T_288 <= _T_287;
    _T_289 <= _T_288;
    _T_290 <= _T_289;
    _T_291 <= _T_290;
    _T_292 <= _T_291;
    _T_293 <= _T_292;
    _T_294 <= _T_293;
    _T_295 <= _T_294;
    _T_296 <= _T_295;
    _T_297 <= _T_296;
    _T_298 <= _T_297;
    _T_299 <= _T_298;
    _T_300 <= io_sig_stat2trans;
    _T_301 <= _T_300;
    _T_302 <= _T_301;
    _T_303 <= _T_302;
    _T_304 <= _T_303;
    _T_305 <= _T_304;
    _T_306 <= _T_305;
    _T_307 <= _T_306;
    _T_308 <= _T_307;
    _T_309 <= _T_308;
    _T_310 <= _T_309;
    _T_311 <= _T_310;
    _T_312 <= _T_311;
    _T_313 <= _T_312;
    _T_314 <= _T_313;
    _T_315 <= io_sig_stat2trans;
    _T_316 <= _T_315;
    _T_317 <= _T_316;
    _T_318 <= _T_317;
    _T_319 <= _T_318;
    _T_320 <= _T_319;
    _T_321 <= _T_320;
    _T_322 <= _T_321;
    _T_323 <= _T_322;
    _T_324 <= _T_323;
    _T_325 <= _T_324;
    _T_326 <= _T_325;
    _T_327 <= _T_326;
    _T_328 <= _T_327;
    _T_329 <= _T_328;
    _T_330 <= io_sig_stat2trans;
    _T_331 <= _T_330;
    _T_332 <= _T_331;
    _T_333 <= _T_332;
    _T_334 <= _T_333;
    _T_335 <= _T_334;
    _T_336 <= _T_335;
    _T_337 <= _T_336;
    _T_338 <= _T_337;
    _T_339 <= _T_338;
    _T_340 <= _T_339;
    _T_341 <= _T_340;
    _T_342 <= _T_341;
    _T_343 <= _T_342;
    _T_344 <= _T_343;
    _T_345 <= io_sig_stat2trans;
    _T_346 <= _T_345;
    _T_347 <= _T_346;
    _T_348 <= _T_347;
    _T_349 <= _T_348;
    _T_350 <= _T_349;
    _T_351 <= _T_350;
    _T_352 <= _T_351;
    _T_353 <= _T_352;
    _T_354 <= _T_353;
    _T_355 <= _T_354;
    _T_356 <= _T_355;
    _T_357 <= _T_356;
    _T_358 <= _T_357;
    _T_359 <= _T_358;
    _T_360 <= io_sig_stat2trans;
    _T_361 <= _T_360;
    _T_362 <= _T_361;
    _T_363 <= _T_362;
    _T_364 <= _T_363;
    _T_365 <= _T_364;
    _T_366 <= _T_365;
    _T_367 <= _T_366;
    _T_368 <= _T_367;
    _T_369 <= _T_368;
    _T_370 <= _T_369;
    _T_371 <= _T_370;
    _T_372 <= _T_371;
    _T_373 <= _T_372;
    _T_374 <= _T_373;
    _T_375 <= io_sig_stat2trans;
    _T_376 <= _T_375;
    _T_377 <= _T_376;
    _T_378 <= _T_377;
    _T_379 <= _T_378;
    _T_380 <= _T_379;
    _T_381 <= _T_380;
    _T_382 <= _T_381;
    _T_383 <= _T_382;
    _T_384 <= _T_383;
    _T_385 <= _T_384;
    _T_386 <= _T_385;
    _T_387 <= _T_386;
    _T_388 <= _T_387;
    _T_389 <= _T_388;
    _T_390 <= io_sig_stat2trans;
    _T_391 <= _T_390;
    _T_392 <= _T_391;
    _T_393 <= _T_392;
    _T_394 <= _T_393;
    _T_395 <= _T_394;
    _T_396 <= _T_395;
    _T_397 <= _T_396;
    _T_398 <= _T_397;
    _T_399 <= _T_398;
    _T_400 <= _T_399;
    _T_401 <= _T_400;
    _T_402 <= _T_401;
    _T_403 <= _T_402;
    _T_404 <= _T_403;
    _T_405 <= io_sig_stat2trans;
    _T_406 <= _T_405;
    _T_407 <= _T_406;
    _T_408 <= _T_407;
    _T_409 <= _T_408;
    _T_410 <= _T_409;
    _T_411 <= _T_410;
    _T_412 <= _T_411;
    _T_413 <= _T_412;
    _T_414 <= _T_413;
    _T_415 <= _T_414;
    _T_416 <= _T_415;
    _T_417 <= _T_416;
    _T_418 <= _T_417;
    _T_419 <= _T_418;
    _T_420 <= io_sig_stat2trans;
    _T_421 <= _T_420;
    _T_422 <= _T_421;
    _T_423 <= _T_422;
    _T_424 <= _T_423;
    _T_425 <= _T_424;
    _T_426 <= _T_425;
    _T_427 <= _T_426;
    _T_428 <= _T_427;
    _T_429 <= _T_428;
    _T_430 <= _T_429;
    _T_431 <= _T_430;
    _T_432 <= _T_431;
    _T_433 <= _T_432;
    _T_434 <= _T_433;
    _T_435 <= io_sig_stat2trans;
    _T_436 <= _T_435;
    _T_437 <= _T_436;
    _T_438 <= _T_437;
    _T_439 <= _T_438;
    _T_440 <= _T_439;
    _T_441 <= _T_440;
    _T_442 <= _T_441;
    _T_443 <= _T_442;
    _T_444 <= _T_443;
    _T_445 <= _T_444;
    _T_446 <= _T_445;
    _T_447 <= _T_446;
    _T_448 <= _T_447;
    _T_449 <= _T_448;
    _T_450 <= io_sig_stat2trans;
    _T_451 <= _T_450;
    _T_452 <= _T_451;
    _T_453 <= _T_452;
    _T_454 <= _T_453;
    _T_455 <= _T_454;
    _T_456 <= _T_455;
    _T_457 <= _T_456;
    _T_458 <= _T_457;
    _T_459 <= _T_458;
    _T_460 <= _T_459;
    _T_461 <= _T_460;
    _T_462 <= _T_461;
    _T_463 <= _T_462;
    _T_464 <= _T_463;
    _T_465 <= io_sig_stat2trans;
    _T_466 <= _T_465;
    _T_467 <= _T_466;
    _T_468 <= _T_467;
    _T_469 <= _T_468;
    _T_470 <= _T_469;
    _T_471 <= _T_470;
    _T_472 <= _T_471;
    _T_473 <= _T_472;
    _T_474 <= _T_473;
    _T_475 <= _T_474;
    _T_476 <= _T_475;
    _T_477 <= _T_476;
    _T_478 <= _T_477;
    _T_479 <= _T_478;
    _T_480 <= io_sig_stat2trans;
    _T_481 <= _T_480;
    _T_482 <= _T_481;
    _T_483 <= _T_482;
    _T_484 <= _T_483;
    _T_485 <= _T_484;
    _T_486 <= _T_485;
    _T_487 <= _T_486;
    _T_488 <= _T_487;
    _T_489 <= _T_488;
    _T_490 <= _T_489;
    _T_491 <= _T_490;
    _T_492 <= _T_491;
    _T_493 <= _T_492;
    _T_494 <= _T_493;
    _T_495 <= io_sig_stat2trans;
    _T_496 <= _T_495;
    _T_497 <= _T_496;
    _T_498 <= _T_497;
    _T_499 <= _T_498;
    _T_500 <= _T_499;
    _T_501 <= _T_500;
    _T_502 <= _T_501;
    _T_503 <= _T_502;
    _T_504 <= _T_503;
    _T_505 <= _T_504;
    _T_506 <= _T_505;
    _T_507 <= _T_506;
    _T_508 <= _T_507;
    _T_509 <= _T_508;
    _T_510 <= io_sig_stat2trans;
    _T_511 <= _T_510;
    _T_512 <= _T_511;
    _T_513 <= _T_512;
    _T_514 <= _T_513;
    _T_515 <= _T_514;
    _T_516 <= _T_515;
    _T_517 <= _T_516;
    _T_518 <= _T_517;
    _T_519 <= _T_518;
    _T_520 <= _T_519;
    _T_521 <= _T_520;
    _T_522 <= _T_521;
    _T_523 <= _T_522;
    _T_524 <= _T_523;
    _T_525 <= io_sig_stat2trans;
    _T_526 <= _T_525;
    _T_527 <= _T_526;
    _T_528 <= _T_527;
    _T_529 <= _T_528;
    _T_530 <= _T_529;
    _T_531 <= _T_530;
    _T_532 <= _T_531;
    _T_533 <= _T_532;
    _T_534 <= _T_533;
    _T_535 <= _T_534;
    _T_536 <= _T_535;
    _T_537 <= _T_536;
    _T_538 <= _T_537;
    _T_539 <= _T_538;
    _T_540 <= io_sig_stat2trans;
    _T_541 <= _T_540;
    _T_542 <= _T_541;
    _T_543 <= _T_542;
    _T_544 <= _T_543;
    _T_545 <= _T_544;
    _T_546 <= _T_545;
    _T_547 <= _T_546;
    _T_548 <= _T_547;
    _T_549 <= _T_548;
    _T_550 <= _T_549;
    _T_551 <= _T_550;
    _T_552 <= _T_551;
    _T_553 <= _T_552;
    _T_554 <= _T_553;
    _T_555 <= io_sig_stat2trans;
    _T_556 <= _T_555;
    _T_557 <= _T_556;
    _T_558 <= _T_557;
    _T_559 <= _T_558;
    _T_560 <= _T_559;
    _T_561 <= _T_560;
    _T_562 <= _T_561;
    _T_563 <= _T_562;
    _T_564 <= _T_563;
    _T_565 <= _T_564;
    _T_566 <= _T_565;
    _T_567 <= _T_566;
    _T_568 <= _T_567;
    _T_569 <= _T_568;
  end
endmodule
module MultiDimMem(
  input         clock,
  input         reset,
  input         io_rd_addr_valid,
  input  [1:0]  io_rd_addr_bits_0,
  input  [1:0]  io_rd_addr_bits_1,
  input  [1:0]  io_rd_addr_bits_2,
  output        io_rd_data_valid,
  output [15:0] io_rd_data_bits,
  input         io_wr_addr_valid,
  input  [1:0]  io_wr_addr_bits_0,
  input  [1:0]  io_wr_addr_bits_1,
  input  [1:0]  io_wr_addr_bits_2,
  input         io_wr_data_valid,
  input  [15:0] io_wr_data_bits
);
  reg [16:0] mem [0:3071]; // @[mem.scala 116:24]
  reg [31:0] _RAND_0;
  wire [16:0] mem_mem_output_data; // @[mem.scala 116:24]
  wire [11:0] mem_mem_output_addr; // @[mem.scala 116:24]
  reg [31:0] _RAND_1;
  wire [16:0] mem__T_61_data; // @[mem.scala 116:24]
  wire [11:0] mem__T_61_addr; // @[mem.scala 116:24]
  wire  mem__T_61_mask; // @[mem.scala 116:24]
  wire  mem__T_61_en; // @[mem.scala 116:24]
  reg  mem_mem_output_en_pipe_0;
  reg [31:0] _RAND_2;
  reg [11:0] mem_mem_output_addr_pipe_0;
  reg [31:0] _RAND_3;
  reg  rd_addr_reg_valid; // @[mem.scala 117:28]
  reg [31:0] _RAND_4;
  reg [15:0] rd_addr_reg_bits_2; // @[mem.scala 117:28]
  reg [31:0] _RAND_5;
  reg [15:0] rd_addr_reg_bits_1; // @[mem.scala 117:28]
  reg [31:0] _RAND_6;
  reg [15:0] rd_addr_reg_bits_0; // @[mem.scala 117:28]
  reg [31:0] _RAND_7;
  wire [15:0] _T_8 = rd_addr_reg_bits_0 + 16'h1; // @[mem.scala 128:102]
  wire  _T_9 = 2'h1 == io_rd_addr_bits_0; // @[Mux.scala 68:19]
  wire  _T_11 = 2'h0 == io_rd_addr_bits_0; // @[Mux.scala 68:19]
  wire [15:0] _T_13 = rd_addr_reg_bits_1 + 16'hc; // @[mem.scala 128:102]
  wire  _T_14 = 2'h1 == io_rd_addr_bits_1; // @[Mux.scala 68:19]
  wire  _T_16 = 2'h0 == io_rd_addr_bits_1; // @[Mux.scala 68:19]
  wire [15:0] _T_18 = rd_addr_reg_bits_2 + 16'hc0; // @[mem.scala 128:102]
  wire  _T_19 = 2'h1 == io_rd_addr_bits_2; // @[Mux.scala 68:19]
  wire  _T_21 = 2'h0 == io_rd_addr_bits_2; // @[Mux.scala 68:19]
  wire [15:0] _T_23 = rd_addr_reg_bits_0 + rd_addr_reg_bits_1; // @[mem.scala 132:46]
  wire [15:0] mem_rd_addr = _T_23 + rd_addr_reg_bits_2; // @[mem.scala 132:46]
  reg  mem_req_valid; // @[mem.scala 139:30]
  reg [31:0] _RAND_8;
  reg  wr_addr_reg_valid; // @[mem.scala 142:28]
  reg [31:0] _RAND_9;
  reg [15:0] wr_addr_reg_bits_2; // @[mem.scala 142:28]
  reg [31:0] _RAND_10;
  reg [15:0] wr_addr_reg_bits_1; // @[mem.scala 142:28]
  reg [31:0] _RAND_11;
  reg [15:0] wr_addr_reg_bits_0; // @[mem.scala 142:28]
  reg [31:0] _RAND_12;
  wire [15:0] _T_40 = wr_addr_reg_bits_0 + 16'h1; // @[mem.scala 154:102]
  wire  _T_41 = 2'h1 == io_wr_addr_bits_0; // @[Mux.scala 68:19]
  wire  _T_43 = 2'h0 == io_wr_addr_bits_0; // @[Mux.scala 68:19]
  wire [15:0] _T_45 = wr_addr_reg_bits_1 + 16'hc; // @[mem.scala 154:102]
  wire  _T_46 = 2'h1 == io_wr_addr_bits_1; // @[Mux.scala 68:19]
  wire  _T_48 = 2'h0 == io_wr_addr_bits_1; // @[Mux.scala 68:19]
  wire [15:0] _T_50 = wr_addr_reg_bits_2 + 16'hc0; // @[mem.scala 154:102]
  wire  _T_51 = 2'h1 == io_wr_addr_bits_2; // @[Mux.scala 68:19]
  wire  _T_53 = 2'h0 == io_wr_addr_bits_2; // @[Mux.scala 68:19]
  reg  wr_data_reg_valid; // @[mem.scala 161:28]
  reg [31:0] _RAND_13;
  reg [15:0] wr_data_reg_bits; // @[mem.scala 161:28]
  reg [31:0] _RAND_14;
  wire [15:0] _T_56 = wr_addr_reg_bits_0 + wr_addr_reg_bits_1; // @[mem.scala 162:46]
  wire [15:0] mem_wr_addr = _T_56 + wr_addr_reg_bits_2; // @[mem.scala 162:46]
  wire [16:0] _GEN_9 = {wr_data_reg_valid, 16'h0}; // @[mem.scala 165:47]
  wire [31:0] _T_58 = {{15'd0}, _GEN_9}; // @[mem.scala 165:47]
  wire [31:0] _GEN_10 = {{16'd0}, wr_data_reg_bits}; // @[mem.scala 165:61]
  wire [31:0] _T_59 = _T_58 | _GEN_10; // @[mem.scala 165:61]
  wire  _T_63 = ~reset; // @[mem.scala 167:9]
  assign mem_mem_output_addr = mem_mem_output_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_mem_output_data = mem[mem_mem_output_addr]; // @[mem.scala 116:24]
  `else
  assign mem_mem_output_data = mem_mem_output_addr >= 12'hc00 ? _RAND_1[16:0] : mem[mem_mem_output_addr]; // @[mem.scala 116:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem__T_61_data = _T_59[16:0];
  assign mem__T_61_addr = mem_wr_addr[11:0];
  assign mem__T_61_mask = 1'h1;
  assign mem__T_61_en = wr_addr_reg_valid;
  assign io_rd_data_valid = mem_req_valid & mem_mem_output_data[16]; // @[mem.scala 140:20]
  assign io_rd_data_bits = mem_req_valid ? mem_mem_output_data[15:0] : 16'h0; // @[mem.scala 141:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3072; initvar = initvar+1)
    mem[initvar] = _RAND_0[16:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  mem_mem_output_en_pipe_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  mem_mem_output_addr_pipe_0 = _RAND_3[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  rd_addr_reg_valid = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  rd_addr_reg_bits_2 = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  rd_addr_reg_bits_1 = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  rd_addr_reg_bits_0 = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  mem_req_valid = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  wr_addr_reg_valid = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  wr_addr_reg_bits_2 = _RAND_10[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  wr_addr_reg_bits_1 = _RAND_11[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  wr_addr_reg_bits_0 = _RAND_12[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  wr_data_reg_valid = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  wr_data_reg_bits = _RAND_14[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(mem__T_61_en & mem__T_61_mask) begin
      mem[mem__T_61_addr] <= mem__T_61_data; // @[mem.scala 116:24]
    end
    mem_mem_output_en_pipe_0 <= rd_addr_reg_valid;
    if (rd_addr_reg_valid) begin
      mem_mem_output_addr_pipe_0 <= mem_rd_addr[11:0];
    end
    if (reset) begin
      rd_addr_reg_valid <= 1'h0;
    end else begin
      rd_addr_reg_valid <= io_rd_addr_valid;
    end
    if (reset) begin
      rd_addr_reg_bits_2 <= 16'h0;
    end else if (_T_21) begin
      rd_addr_reg_bits_2 <= 16'h0;
    end else if (_T_19) begin
      rd_addr_reg_bits_2 <= _T_18;
    end
    if (reset) begin
      rd_addr_reg_bits_1 <= 16'h0;
    end else if (_T_16) begin
      rd_addr_reg_bits_1 <= 16'h0;
    end else if (_T_14) begin
      rd_addr_reg_bits_1 <= _T_13;
    end
    if (reset) begin
      rd_addr_reg_bits_0 <= 16'h0;
    end else if (_T_11) begin
      rd_addr_reg_bits_0 <= 16'h0;
    end else if (_T_9) begin
      rd_addr_reg_bits_0 <= _T_8;
    end
    if (reset) begin
      mem_req_valid <= 1'h0;
    end else begin
      mem_req_valid <= rd_addr_reg_valid;
    end
    if (reset) begin
      wr_addr_reg_valid <= 1'h0;
    end else begin
      wr_addr_reg_valid <= io_wr_addr_valid;
    end
    if (reset) begin
      wr_addr_reg_bits_2 <= 16'h0;
    end else if (_T_53) begin
      wr_addr_reg_bits_2 <= 16'h0;
    end else if (_T_51) begin
      wr_addr_reg_bits_2 <= _T_50;
    end
    if (reset) begin
      wr_addr_reg_bits_1 <= 16'h0;
    end else if (_T_48) begin
      wr_addr_reg_bits_1 <= 16'h0;
    end else if (_T_46) begin
      wr_addr_reg_bits_1 <= _T_45;
    end
    if (reset) begin
      wr_addr_reg_bits_0 <= 16'h0;
    end else if (_T_43) begin
      wr_addr_reg_bits_0 <= 16'h0;
    end else if (_T_41) begin
      wr_addr_reg_bits_0 <= _T_40;
    end
    if (reset) begin
      wr_data_reg_valid <= 1'h0;
    end else begin
      wr_data_reg_valid <= io_wr_data_valid;
    end
    if (reset) begin
      wr_data_reg_bits <= 16'h0;
    end else begin
      wr_data_reg_bits <= io_wr_data_bits;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_63) begin
          $fwrite(32'h80000002,"wr_addr:%d %d, wr_data: %d, rd_addr:%d %d, rd_data: %d %d\n",mem_wr_addr,wr_addr_reg_valid,wr_data_reg_bits,mem_rd_addr,rd_addr_reg_valid,io_rd_data_valid,io_rd_data_bits); // @[mem.scala 167:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module MemController(
  input         clock,
  input         reset,
  input         io_rd_valid,
  input         io_wr_valid,
  output        io_rd_data_valid,
  output [15:0] io_rd_data_bits,
  input         io_wr_data_valid,
  input  [15:0] io_wr_data_bits
);
  wire  MultiDimMem_clock; // @[mem.scala 31:19]
  wire  MultiDimMem_reset; // @[mem.scala 31:19]
  wire  MultiDimMem_io_rd_addr_valid; // @[mem.scala 31:19]
  wire [1:0] MultiDimMem_io_rd_addr_bits_0; // @[mem.scala 31:19]
  wire [1:0] MultiDimMem_io_rd_addr_bits_1; // @[mem.scala 31:19]
  wire [1:0] MultiDimMem_io_rd_addr_bits_2; // @[mem.scala 31:19]
  wire  MultiDimMem_io_rd_data_valid; // @[mem.scala 31:19]
  wire [15:0] MultiDimMem_io_rd_data_bits; // @[mem.scala 31:19]
  wire  MultiDimMem_io_wr_addr_valid; // @[mem.scala 31:19]
  wire [1:0] MultiDimMem_io_wr_addr_bits_0; // @[mem.scala 31:19]
  wire [1:0] MultiDimMem_io_wr_addr_bits_1; // @[mem.scala 31:19]
  wire [1:0] MultiDimMem_io_wr_addr_bits_2; // @[mem.scala 31:19]
  wire  MultiDimMem_io_wr_data_valid; // @[mem.scala 31:19]
  wire [15:0] MultiDimMem_io_wr_data_bits; // @[mem.scala 31:19]
  wire  MultiDimTime_clock; // @[mem.scala 32:23]
  wire  MultiDimTime_reset; // @[mem.scala 32:23]
  wire  MultiDimTime_io_in; // @[mem.scala 32:23]
  wire [1:0] MultiDimTime_io_out_0; // @[mem.scala 32:23]
  wire [1:0] MultiDimTime_io_out_1; // @[mem.scala 32:23]
  wire [1:0] MultiDimTime_io_out_2; // @[mem.scala 32:23]
  wire [15:0] MultiDimTime_io_index_0; // @[mem.scala 32:23]
  wire [15:0] MultiDimTime_io_index_1; // @[mem.scala 32:23]
  wire [15:0] MultiDimTime_io_index_2; // @[mem.scala 32:23]
  wire  MultiDimTime_1_clock; // @[mem.scala 33:23]
  wire  MultiDimTime_1_reset; // @[mem.scala 33:23]
  wire  MultiDimTime_1_io_in; // @[mem.scala 33:23]
  wire [1:0] MultiDimTime_1_io_out_0; // @[mem.scala 33:23]
  wire [1:0] MultiDimTime_1_io_out_1; // @[mem.scala 33:23]
  wire [1:0] MultiDimTime_1_io_out_2; // @[mem.scala 33:23]
  wire [15:0] MultiDimTime_1_io_index_0; // @[mem.scala 33:23]
  wire [15:0] MultiDimTime_1_io_index_1; // @[mem.scala 33:23]
  wire [15:0] MultiDimTime_1_io_index_2; // @[mem.scala 33:23]
  MultiDimMem MultiDimMem ( // @[mem.scala 31:19]
    .clock(MultiDimMem_clock),
    .reset(MultiDimMem_reset),
    .io_rd_addr_valid(MultiDimMem_io_rd_addr_valid),
    .io_rd_addr_bits_0(MultiDimMem_io_rd_addr_bits_0),
    .io_rd_addr_bits_1(MultiDimMem_io_rd_addr_bits_1),
    .io_rd_addr_bits_2(MultiDimMem_io_rd_addr_bits_2),
    .io_rd_data_valid(MultiDimMem_io_rd_data_valid),
    .io_rd_data_bits(MultiDimMem_io_rd_data_bits),
    .io_wr_addr_valid(MultiDimMem_io_wr_addr_valid),
    .io_wr_addr_bits_0(MultiDimMem_io_wr_addr_bits_0),
    .io_wr_addr_bits_1(MultiDimMem_io_wr_addr_bits_1),
    .io_wr_addr_bits_2(MultiDimMem_io_wr_addr_bits_2),
    .io_wr_data_valid(MultiDimMem_io_wr_data_valid),
    .io_wr_data_bits(MultiDimMem_io_wr_data_bits)
  );
  MultiDimTime MultiDimTime ( // @[mem.scala 32:23]
    .clock(MultiDimTime_clock),
    .reset(MultiDimTime_reset),
    .io_in(MultiDimTime_io_in),
    .io_out_0(MultiDimTime_io_out_0),
    .io_out_1(MultiDimTime_io_out_1),
    .io_out_2(MultiDimTime_io_out_2),
    .io_index_0(MultiDimTime_io_index_0),
    .io_index_1(MultiDimTime_io_index_1),
    .io_index_2(MultiDimTime_io_index_2)
  );
  MultiDimTime MultiDimTime_1 ( // @[mem.scala 33:23]
    .clock(MultiDimTime_1_clock),
    .reset(MultiDimTime_1_reset),
    .io_in(MultiDimTime_1_io_in),
    .io_out_0(MultiDimTime_1_io_out_0),
    .io_out_1(MultiDimTime_1_io_out_1),
    .io_out_2(MultiDimTime_1_io_out_2),
    .io_index_0(MultiDimTime_1_io_index_0),
    .io_index_1(MultiDimTime_1_io_index_1),
    .io_index_2(MultiDimTime_1_io_index_2)
  );
  assign io_rd_data_valid = MultiDimMem_io_rd_data_valid; // @[mem.scala 50:14]
  assign io_rd_data_bits = MultiDimMem_io_rd_data_bits; // @[mem.scala 50:14]
  assign MultiDimMem_clock = clock;
  assign MultiDimMem_reset = reset;
  assign MultiDimMem_io_rd_addr_valid = io_rd_valid; // @[mem.scala 47:21]
  assign MultiDimMem_io_rd_addr_bits_0 = MultiDimTime_1_io_out_0; // @[mem.scala 46:20]
  assign MultiDimMem_io_rd_addr_bits_1 = MultiDimTime_1_io_out_1; // @[mem.scala 46:20]
  assign MultiDimMem_io_rd_addr_bits_2 = MultiDimTime_1_io_out_2; // @[mem.scala 46:20]
  assign MultiDimMem_io_wr_addr_valid = io_wr_valid; // @[mem.scala 43:21]
  assign MultiDimMem_io_wr_addr_bits_0 = MultiDimTime_io_out_0; // @[mem.scala 42:20]
  assign MultiDimMem_io_wr_addr_bits_1 = MultiDimTime_io_out_1; // @[mem.scala 42:20]
  assign MultiDimMem_io_wr_addr_bits_2 = MultiDimTime_io_out_2; // @[mem.scala 42:20]
  assign MultiDimMem_io_wr_data_valid = io_wr_data_valid; // @[mem.scala 51:15]
  assign MultiDimMem_io_wr_data_bits = io_wr_data_bits; // @[mem.scala 51:15]
  assign MultiDimTime_clock = clock;
  assign MultiDimTime_reset = reset;
  assign MultiDimTime_io_in = io_wr_valid; // @[mem.scala 41:14]
  assign MultiDimTime_1_clock = clock;
  assign MultiDimTime_1_reset = reset;
  assign MultiDimTime_1_io_in = io_rd_valid; // @[mem.scala 45:14]
endmodule
module MultiDimMem_22(
  input          clock,
  input          reset,
  input          io_rd_addr_valid,
  input  [1:0]   io_rd_addr_bits_0,
  input  [1:0]   io_rd_addr_bits_1,
  input  [1:0]   io_rd_addr_bits_2,
  output         io_rd_data_valid,
  output [127:0] io_rd_data_bits,
  input          io_wr_addr_valid,
  input  [1:0]   io_wr_addr_bits_0,
  input  [1:0]   io_wr_addr_bits_1,
  input  [1:0]   io_wr_addr_bits_2,
  input          io_wr_data_valid,
  input  [127:0] io_wr_data_bits
);
  reg [128:0] mem [0:3071]; // @[mem.scala 116:24]
  reg [159:0] _RAND_0;
  wire [128:0] mem_mem_output_data; // @[mem.scala 116:24]
  wire [11:0] mem_mem_output_addr; // @[mem.scala 116:24]
  reg [159:0] _RAND_1;
  wire [128:0] mem__T_61_data; // @[mem.scala 116:24]
  wire [11:0] mem__T_61_addr; // @[mem.scala 116:24]
  wire  mem__T_61_mask; // @[mem.scala 116:24]
  wire  mem__T_61_en; // @[mem.scala 116:24]
  reg  mem_mem_output_en_pipe_0;
  reg [31:0] _RAND_2;
  reg [11:0] mem_mem_output_addr_pipe_0;
  reg [31:0] _RAND_3;
  reg  rd_addr_reg_valid; // @[mem.scala 117:28]
  reg [31:0] _RAND_4;
  reg [15:0] rd_addr_reg_bits_2; // @[mem.scala 117:28]
  reg [31:0] _RAND_5;
  reg [15:0] rd_addr_reg_bits_1; // @[mem.scala 117:28]
  reg [31:0] _RAND_6;
  reg [15:0] rd_addr_reg_bits_0; // @[mem.scala 117:28]
  reg [31:0] _RAND_7;
  wire [15:0] _T_8 = rd_addr_reg_bits_0 + 16'h1; // @[mem.scala 128:102]
  wire  _T_9 = 2'h1 == io_rd_addr_bits_0; // @[Mux.scala 68:19]
  wire  _T_11 = 2'h0 == io_rd_addr_bits_0; // @[Mux.scala 68:19]
  wire [15:0] _T_13 = rd_addr_reg_bits_1 + 16'hc; // @[mem.scala 128:102]
  wire  _T_14 = 2'h1 == io_rd_addr_bits_1; // @[Mux.scala 68:19]
  wire  _T_16 = 2'h0 == io_rd_addr_bits_1; // @[Mux.scala 68:19]
  wire [15:0] _T_18 = rd_addr_reg_bits_2 + 16'hc0; // @[mem.scala 128:102]
  wire  _T_19 = 2'h1 == io_rd_addr_bits_2; // @[Mux.scala 68:19]
  wire  _T_21 = 2'h0 == io_rd_addr_bits_2; // @[Mux.scala 68:19]
  wire [15:0] _T_23 = rd_addr_reg_bits_0 + rd_addr_reg_bits_1; // @[mem.scala 132:46]
  wire [15:0] mem_rd_addr = _T_23 + rd_addr_reg_bits_2; // @[mem.scala 132:46]
  reg  mem_req_valid; // @[mem.scala 139:30]
  reg [31:0] _RAND_8;
  reg  wr_addr_reg_valid; // @[mem.scala 142:28]
  reg [31:0] _RAND_9;
  reg [15:0] wr_addr_reg_bits_2; // @[mem.scala 142:28]
  reg [31:0] _RAND_10;
  reg [15:0] wr_addr_reg_bits_1; // @[mem.scala 142:28]
  reg [31:0] _RAND_11;
  reg [15:0] wr_addr_reg_bits_0; // @[mem.scala 142:28]
  reg [31:0] _RAND_12;
  wire [15:0] _T_40 = wr_addr_reg_bits_0 + 16'h1; // @[mem.scala 154:102]
  wire  _T_41 = 2'h1 == io_wr_addr_bits_0; // @[Mux.scala 68:19]
  wire  _T_43 = 2'h0 == io_wr_addr_bits_0; // @[Mux.scala 68:19]
  wire [15:0] _T_45 = wr_addr_reg_bits_1 + 16'hc; // @[mem.scala 154:102]
  wire  _T_46 = 2'h1 == io_wr_addr_bits_1; // @[Mux.scala 68:19]
  wire  _T_48 = 2'h0 == io_wr_addr_bits_1; // @[Mux.scala 68:19]
  wire [15:0] _T_50 = wr_addr_reg_bits_2 + 16'hc0; // @[mem.scala 154:102]
  wire  _T_51 = 2'h1 == io_wr_addr_bits_2; // @[Mux.scala 68:19]
  wire  _T_53 = 2'h0 == io_wr_addr_bits_2; // @[Mux.scala 68:19]
  reg  wr_data_reg_valid; // @[mem.scala 161:28]
  reg [31:0] _RAND_13;
  reg [127:0] wr_data_reg_bits; // @[mem.scala 161:28]
  reg [127:0] _RAND_14;
  wire [15:0] _T_56 = wr_addr_reg_bits_0 + wr_addr_reg_bits_1; // @[mem.scala 162:46]
  wire [15:0] mem_wr_addr = _T_56 + wr_addr_reg_bits_2; // @[mem.scala 162:46]
  wire [128:0] _GEN_9 = {wr_data_reg_valid, 128'h0}; // @[mem.scala 165:47]
  wire [255:0] _T_58 = {{127'd0}, _GEN_9}; // @[mem.scala 165:47]
  wire [255:0] _GEN_10 = {{128'd0}, wr_data_reg_bits}; // @[mem.scala 165:61]
  wire [255:0] _T_59 = _T_58 | _GEN_10; // @[mem.scala 165:61]
  wire  _T_63 = ~reset; // @[mem.scala 167:9]
  assign mem_mem_output_addr = mem_mem_output_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_mem_output_data = mem[mem_mem_output_addr]; // @[mem.scala 116:24]
  `else
  assign mem_mem_output_data = mem_mem_output_addr >= 12'hc00 ? _RAND_1[128:0] : mem[mem_mem_output_addr]; // @[mem.scala 116:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem__T_61_data = _T_59[128:0];
  assign mem__T_61_addr = mem_wr_addr[11:0];
  assign mem__T_61_mask = 1'h1;
  assign mem__T_61_en = wr_addr_reg_valid;
  assign io_rd_data_valid = mem_req_valid & mem_mem_output_data[128]; // @[mem.scala 140:20]
  assign io_rd_data_bits = mem_req_valid ? mem_mem_output_data[127:0] : 128'h0; // @[mem.scala 141:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {5{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3072; initvar = initvar+1)
    mem[initvar] = _RAND_0[128:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {5{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  mem_mem_output_en_pipe_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  mem_mem_output_addr_pipe_0 = _RAND_3[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  rd_addr_reg_valid = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  rd_addr_reg_bits_2 = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  rd_addr_reg_bits_1 = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  rd_addr_reg_bits_0 = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  mem_req_valid = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  wr_addr_reg_valid = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  wr_addr_reg_bits_2 = _RAND_10[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  wr_addr_reg_bits_1 = _RAND_11[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  wr_addr_reg_bits_0 = _RAND_12[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  wr_data_reg_valid = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {4{`RANDOM}};
  wr_data_reg_bits = _RAND_14[127:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(mem__T_61_en & mem__T_61_mask) begin
      mem[mem__T_61_addr] <= mem__T_61_data; // @[mem.scala 116:24]
    end
    mem_mem_output_en_pipe_0 <= rd_addr_reg_valid;
    if (rd_addr_reg_valid) begin
      mem_mem_output_addr_pipe_0 <= mem_rd_addr[11:0];
    end
    if (reset) begin
      rd_addr_reg_valid <= 1'h0;
    end else begin
      rd_addr_reg_valid <= io_rd_addr_valid;
    end
    if (reset) begin
      rd_addr_reg_bits_2 <= 16'h0;
    end else if (_T_21) begin
      rd_addr_reg_bits_2 <= 16'h0;
    end else if (_T_19) begin
      rd_addr_reg_bits_2 <= _T_18;
    end
    if (reset) begin
      rd_addr_reg_bits_1 <= 16'h0;
    end else if (_T_16) begin
      rd_addr_reg_bits_1 <= 16'h0;
    end else if (_T_14) begin
      rd_addr_reg_bits_1 <= _T_13;
    end
    if (reset) begin
      rd_addr_reg_bits_0 <= 16'h0;
    end else if (_T_11) begin
      rd_addr_reg_bits_0 <= 16'h0;
    end else if (_T_9) begin
      rd_addr_reg_bits_0 <= _T_8;
    end
    if (reset) begin
      mem_req_valid <= 1'h0;
    end else begin
      mem_req_valid <= rd_addr_reg_valid;
    end
    if (reset) begin
      wr_addr_reg_valid <= 1'h0;
    end else begin
      wr_addr_reg_valid <= io_wr_addr_valid;
    end
    if (reset) begin
      wr_addr_reg_bits_2 <= 16'h0;
    end else if (_T_53) begin
      wr_addr_reg_bits_2 <= 16'h0;
    end else if (_T_51) begin
      wr_addr_reg_bits_2 <= _T_50;
    end
    if (reset) begin
      wr_addr_reg_bits_1 <= 16'h0;
    end else if (_T_48) begin
      wr_addr_reg_bits_1 <= 16'h0;
    end else if (_T_46) begin
      wr_addr_reg_bits_1 <= _T_45;
    end
    if (reset) begin
      wr_addr_reg_bits_0 <= 16'h0;
    end else if (_T_43) begin
      wr_addr_reg_bits_0 <= 16'h0;
    end else if (_T_41) begin
      wr_addr_reg_bits_0 <= _T_40;
    end
    if (reset) begin
      wr_data_reg_valid <= 1'h0;
    end else begin
      wr_data_reg_valid <= io_wr_data_valid;
    end
    if (reset) begin
      wr_data_reg_bits <= 128'h0;
    end else begin
      wr_data_reg_bits <= io_wr_data_bits;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_63) begin
          $fwrite(32'h80000002,"wr_addr:%d %d, wr_data: %d, rd_addr:%d %d, rd_data: %d %d\n",mem_wr_addr,wr_addr_reg_valid,wr_data_reg_bits,mem_rd_addr,rd_addr_reg_valid,io_rd_data_valid,io_rd_data_bits); // @[mem.scala 167:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module MemController_22(
  input          clock,
  input          reset,
  input          io_rd_valid,
  input          io_wr_valid,
  output         io_rd_data_valid,
  output [127:0] io_rd_data_bits,
  input          io_wr_data_valid,
  input  [127:0] io_wr_data_bits
);
  wire  MultiDimMem_clock; // @[mem.scala 31:19]
  wire  MultiDimMem_reset; // @[mem.scala 31:19]
  wire  MultiDimMem_io_rd_addr_valid; // @[mem.scala 31:19]
  wire [1:0] MultiDimMem_io_rd_addr_bits_0; // @[mem.scala 31:19]
  wire [1:0] MultiDimMem_io_rd_addr_bits_1; // @[mem.scala 31:19]
  wire [1:0] MultiDimMem_io_rd_addr_bits_2; // @[mem.scala 31:19]
  wire  MultiDimMem_io_rd_data_valid; // @[mem.scala 31:19]
  wire [127:0] MultiDimMem_io_rd_data_bits; // @[mem.scala 31:19]
  wire  MultiDimMem_io_wr_addr_valid; // @[mem.scala 31:19]
  wire [1:0] MultiDimMem_io_wr_addr_bits_0; // @[mem.scala 31:19]
  wire [1:0] MultiDimMem_io_wr_addr_bits_1; // @[mem.scala 31:19]
  wire [1:0] MultiDimMem_io_wr_addr_bits_2; // @[mem.scala 31:19]
  wire  MultiDimMem_io_wr_data_valid; // @[mem.scala 31:19]
  wire [127:0] MultiDimMem_io_wr_data_bits; // @[mem.scala 31:19]
  wire  MultiDimTime_clock; // @[mem.scala 32:23]
  wire  MultiDimTime_reset; // @[mem.scala 32:23]
  wire  MultiDimTime_io_in; // @[mem.scala 32:23]
  wire [1:0] MultiDimTime_io_out_0; // @[mem.scala 32:23]
  wire [1:0] MultiDimTime_io_out_1; // @[mem.scala 32:23]
  wire [1:0] MultiDimTime_io_out_2; // @[mem.scala 32:23]
  wire [15:0] MultiDimTime_io_index_0; // @[mem.scala 32:23]
  wire [15:0] MultiDimTime_io_index_1; // @[mem.scala 32:23]
  wire [15:0] MultiDimTime_io_index_2; // @[mem.scala 32:23]
  wire  MultiDimTime_1_clock; // @[mem.scala 33:23]
  wire  MultiDimTime_1_reset; // @[mem.scala 33:23]
  wire  MultiDimTime_1_io_in; // @[mem.scala 33:23]
  wire [1:0] MultiDimTime_1_io_out_0; // @[mem.scala 33:23]
  wire [1:0] MultiDimTime_1_io_out_1; // @[mem.scala 33:23]
  wire [1:0] MultiDimTime_1_io_out_2; // @[mem.scala 33:23]
  wire [15:0] MultiDimTime_1_io_index_0; // @[mem.scala 33:23]
  wire [15:0] MultiDimTime_1_io_index_1; // @[mem.scala 33:23]
  wire [15:0] MultiDimTime_1_io_index_2; // @[mem.scala 33:23]
  MultiDimMem_22 MultiDimMem ( // @[mem.scala 31:19]
    .clock(MultiDimMem_clock),
    .reset(MultiDimMem_reset),
    .io_rd_addr_valid(MultiDimMem_io_rd_addr_valid),
    .io_rd_addr_bits_0(MultiDimMem_io_rd_addr_bits_0),
    .io_rd_addr_bits_1(MultiDimMem_io_rd_addr_bits_1),
    .io_rd_addr_bits_2(MultiDimMem_io_rd_addr_bits_2),
    .io_rd_data_valid(MultiDimMem_io_rd_data_valid),
    .io_rd_data_bits(MultiDimMem_io_rd_data_bits),
    .io_wr_addr_valid(MultiDimMem_io_wr_addr_valid),
    .io_wr_addr_bits_0(MultiDimMem_io_wr_addr_bits_0),
    .io_wr_addr_bits_1(MultiDimMem_io_wr_addr_bits_1),
    .io_wr_addr_bits_2(MultiDimMem_io_wr_addr_bits_2),
    .io_wr_data_valid(MultiDimMem_io_wr_data_valid),
    .io_wr_data_bits(MultiDimMem_io_wr_data_bits)
  );
  MultiDimTime MultiDimTime ( // @[mem.scala 32:23]
    .clock(MultiDimTime_clock),
    .reset(MultiDimTime_reset),
    .io_in(MultiDimTime_io_in),
    .io_out_0(MultiDimTime_io_out_0),
    .io_out_1(MultiDimTime_io_out_1),
    .io_out_2(MultiDimTime_io_out_2),
    .io_index_0(MultiDimTime_io_index_0),
    .io_index_1(MultiDimTime_io_index_1),
    .io_index_2(MultiDimTime_io_index_2)
  );
  MultiDimTime MultiDimTime_1 ( // @[mem.scala 33:23]
    .clock(MultiDimTime_1_clock),
    .reset(MultiDimTime_1_reset),
    .io_in(MultiDimTime_1_io_in),
    .io_out_0(MultiDimTime_1_io_out_0),
    .io_out_1(MultiDimTime_1_io_out_1),
    .io_out_2(MultiDimTime_1_io_out_2),
    .io_index_0(MultiDimTime_1_io_index_0),
    .io_index_1(MultiDimTime_1_io_index_1),
    .io_index_2(MultiDimTime_1_io_index_2)
  );
  assign io_rd_data_valid = MultiDimMem_io_rd_data_valid; // @[mem.scala 50:14]
  assign io_rd_data_bits = MultiDimMem_io_rd_data_bits; // @[mem.scala 50:14]
  assign MultiDimMem_clock = clock;
  assign MultiDimMem_reset = reset;
  assign MultiDimMem_io_rd_addr_valid = io_rd_valid; // @[mem.scala 47:21]
  assign MultiDimMem_io_rd_addr_bits_0 = MultiDimTime_1_io_out_0; // @[mem.scala 46:20]
  assign MultiDimMem_io_rd_addr_bits_1 = MultiDimTime_1_io_out_1; // @[mem.scala 46:20]
  assign MultiDimMem_io_rd_addr_bits_2 = MultiDimTime_1_io_out_2; // @[mem.scala 46:20]
  assign MultiDimMem_io_wr_addr_valid = io_wr_valid; // @[mem.scala 43:21]
  assign MultiDimMem_io_wr_addr_bits_0 = MultiDimTime_io_out_0; // @[mem.scala 42:20]
  assign MultiDimMem_io_wr_addr_bits_1 = MultiDimTime_io_out_1; // @[mem.scala 42:20]
  assign MultiDimMem_io_wr_addr_bits_2 = MultiDimTime_io_out_2; // @[mem.scala 42:20]
  assign MultiDimMem_io_wr_data_valid = io_wr_data_valid; // @[mem.scala 51:15]
  assign MultiDimMem_io_wr_data_bits = io_wr_data_bits; // @[mem.scala 51:15]
  assign MultiDimTime_clock = clock;
  assign MultiDimTime_reset = reset;
  assign MultiDimTime_io_in = io_wr_valid; // @[mem.scala 41:14]
  assign MultiDimTime_1_clock = clock;
  assign MultiDimTime_1_reset = reset;
  assign MultiDimTime_1_io_in = io_rd_valid; // @[mem.scala 45:14]
endmodule
module MultiDimMem_52(
  input          clock,
  input          reset,
  input          io_rd_addr_valid,
  input  [1:0]   io_rd_addr_bits_0,
  input  [1:0]   io_rd_addr_bits_1,
  input  [1:0]   io_rd_addr_bits_2,
  output         io_rd_data_valid,
  output [127:0] io_rd_data_bits,
  input          io_wr_addr_valid,
  input  [1:0]   io_wr_addr_bits_0,
  input  [1:0]   io_wr_addr_bits_1,
  input  [1:0]   io_wr_addr_bits_2,
  input          io_wr_data_valid,
  input  [127:0] io_wr_data_bits
);
  reg [128:0] mem [0:4223]; // @[mem.scala 116:24]
  reg [159:0] _RAND_0;
  wire [128:0] mem_mem_output_data; // @[mem.scala 116:24]
  wire [12:0] mem_mem_output_addr; // @[mem.scala 116:24]
  reg [159:0] _RAND_1;
  wire [128:0] mem__T_61_data; // @[mem.scala 116:24]
  wire [12:0] mem__T_61_addr; // @[mem.scala 116:24]
  wire  mem__T_61_mask; // @[mem.scala 116:24]
  wire  mem__T_61_en; // @[mem.scala 116:24]
  reg  mem_mem_output_en_pipe_0;
  reg [31:0] _RAND_2;
  reg [12:0] mem_mem_output_addr_pipe_0;
  reg [31:0] _RAND_3;
  reg  rd_addr_reg_valid; // @[mem.scala 117:28]
  reg [31:0] _RAND_4;
  reg [15:0] rd_addr_reg_bits_2; // @[mem.scala 117:28]
  reg [31:0] _RAND_5;
  reg [15:0] rd_addr_reg_bits_1; // @[mem.scala 117:28]
  reg [31:0] _RAND_6;
  reg [15:0] rd_addr_reg_bits_0; // @[mem.scala 117:28]
  reg [31:0] _RAND_7;
  wire [15:0] _T_8 = rd_addr_reg_bits_0 + 16'h1; // @[mem.scala 128:102]
  wire  _T_9 = 2'h1 == io_rd_addr_bits_0; // @[Mux.scala 68:19]
  wire  _T_11 = 2'h0 == io_rd_addr_bits_0; // @[Mux.scala 68:19]
  wire [15:0] _T_13 = rd_addr_reg_bits_1 + 16'hc; // @[mem.scala 128:102]
  wire  _T_14 = 2'h1 == io_rd_addr_bits_1; // @[Mux.scala 68:19]
  wire  _T_16 = 2'h0 == io_rd_addr_bits_1; // @[Mux.scala 68:19]
  wire [15:0] _T_18 = rd_addr_reg_bits_2 + 16'h108; // @[mem.scala 128:102]
  wire  _T_19 = 2'h1 == io_rd_addr_bits_2; // @[Mux.scala 68:19]
  wire  _T_21 = 2'h0 == io_rd_addr_bits_2; // @[Mux.scala 68:19]
  wire [15:0] _T_23 = rd_addr_reg_bits_0 + rd_addr_reg_bits_1; // @[mem.scala 132:46]
  wire [15:0] mem_rd_addr = _T_23 + rd_addr_reg_bits_2; // @[mem.scala 132:46]
  reg  mem_req_valid; // @[mem.scala 139:30]
  reg [31:0] _RAND_8;
  reg  wr_addr_reg_valid; // @[mem.scala 142:28]
  reg [31:0] _RAND_9;
  reg [15:0] wr_addr_reg_bits_2; // @[mem.scala 142:28]
  reg [31:0] _RAND_10;
  reg [15:0] wr_addr_reg_bits_1; // @[mem.scala 142:28]
  reg [31:0] _RAND_11;
  reg [15:0] wr_addr_reg_bits_0; // @[mem.scala 142:28]
  reg [31:0] _RAND_12;
  wire [15:0] _T_40 = wr_addr_reg_bits_0 + 16'h1; // @[mem.scala 154:102]
  wire  _T_41 = 2'h1 == io_wr_addr_bits_0; // @[Mux.scala 68:19]
  wire  _T_43 = 2'h0 == io_wr_addr_bits_0; // @[Mux.scala 68:19]
  wire [15:0] _T_45 = wr_addr_reg_bits_1 + 16'hc; // @[mem.scala 154:102]
  wire  _T_46 = 2'h1 == io_wr_addr_bits_1; // @[Mux.scala 68:19]
  wire  _T_48 = 2'h0 == io_wr_addr_bits_1; // @[Mux.scala 68:19]
  wire [15:0] _T_50 = wr_addr_reg_bits_2 + 16'h108; // @[mem.scala 154:102]
  wire  _T_51 = 2'h1 == io_wr_addr_bits_2; // @[Mux.scala 68:19]
  wire  _T_53 = 2'h0 == io_wr_addr_bits_2; // @[Mux.scala 68:19]
  reg  wr_data_reg_valid; // @[mem.scala 161:28]
  reg [31:0] _RAND_13;
  reg [127:0] wr_data_reg_bits; // @[mem.scala 161:28]
  reg [127:0] _RAND_14;
  wire [15:0] _T_56 = wr_addr_reg_bits_0 + wr_addr_reg_bits_1; // @[mem.scala 162:46]
  wire [15:0] mem_wr_addr = _T_56 + wr_addr_reg_bits_2; // @[mem.scala 162:46]
  wire [128:0] _GEN_9 = {wr_data_reg_valid, 128'h0}; // @[mem.scala 165:47]
  wire [255:0] _T_58 = {{127'd0}, _GEN_9}; // @[mem.scala 165:47]
  wire [255:0] _GEN_10 = {{128'd0}, wr_data_reg_bits}; // @[mem.scala 165:61]
  wire [255:0] _T_59 = _T_58 | _GEN_10; // @[mem.scala 165:61]
  wire  _T_63 = ~reset; // @[mem.scala 167:9]
  assign mem_mem_output_addr = mem_mem_output_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_mem_output_data = mem[mem_mem_output_addr]; // @[mem.scala 116:24]
  `else
  assign mem_mem_output_data = mem_mem_output_addr >= 13'h1080 ? _RAND_1[128:0] : mem[mem_mem_output_addr]; // @[mem.scala 116:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem__T_61_data = _T_59[128:0];
  assign mem__T_61_addr = mem_wr_addr[12:0];
  assign mem__T_61_mask = 1'h1;
  assign mem__T_61_en = wr_addr_reg_valid;
  assign io_rd_data_valid = mem_req_valid & mem_mem_output_data[128]; // @[mem.scala 140:20]
  assign io_rd_data_bits = mem_req_valid ? mem_mem_output_data[127:0] : 128'h0; // @[mem.scala 141:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {5{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 4224; initvar = initvar+1)
    mem[initvar] = _RAND_0[128:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {5{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  mem_mem_output_en_pipe_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  mem_mem_output_addr_pipe_0 = _RAND_3[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  rd_addr_reg_valid = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  rd_addr_reg_bits_2 = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  rd_addr_reg_bits_1 = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  rd_addr_reg_bits_0 = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  mem_req_valid = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  wr_addr_reg_valid = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  wr_addr_reg_bits_2 = _RAND_10[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  wr_addr_reg_bits_1 = _RAND_11[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  wr_addr_reg_bits_0 = _RAND_12[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  wr_data_reg_valid = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {4{`RANDOM}};
  wr_data_reg_bits = _RAND_14[127:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(mem__T_61_en & mem__T_61_mask) begin
      mem[mem__T_61_addr] <= mem__T_61_data; // @[mem.scala 116:24]
    end
    mem_mem_output_en_pipe_0 <= rd_addr_reg_valid;
    if (rd_addr_reg_valid) begin
      mem_mem_output_addr_pipe_0 <= mem_rd_addr[12:0];
    end
    if (reset) begin
      rd_addr_reg_valid <= 1'h0;
    end else begin
      rd_addr_reg_valid <= io_rd_addr_valid;
    end
    if (reset) begin
      rd_addr_reg_bits_2 <= 16'h0;
    end else if (_T_21) begin
      rd_addr_reg_bits_2 <= 16'h0;
    end else if (_T_19) begin
      rd_addr_reg_bits_2 <= _T_18;
    end
    if (reset) begin
      rd_addr_reg_bits_1 <= 16'h0;
    end else if (_T_16) begin
      rd_addr_reg_bits_1 <= 16'h0;
    end else if (_T_14) begin
      rd_addr_reg_bits_1 <= _T_13;
    end
    if (reset) begin
      rd_addr_reg_bits_0 <= 16'h0;
    end else if (_T_11) begin
      rd_addr_reg_bits_0 <= 16'h0;
    end else if (_T_9) begin
      rd_addr_reg_bits_0 <= _T_8;
    end
    if (reset) begin
      mem_req_valid <= 1'h0;
    end else begin
      mem_req_valid <= rd_addr_reg_valid;
    end
    if (reset) begin
      wr_addr_reg_valid <= 1'h0;
    end else begin
      wr_addr_reg_valid <= io_wr_addr_valid;
    end
    if (reset) begin
      wr_addr_reg_bits_2 <= 16'h0;
    end else if (_T_53) begin
      wr_addr_reg_bits_2 <= 16'h0;
    end else if (_T_51) begin
      wr_addr_reg_bits_2 <= _T_50;
    end
    if (reset) begin
      wr_addr_reg_bits_1 <= 16'h0;
    end else if (_T_48) begin
      wr_addr_reg_bits_1 <= 16'h0;
    end else if (_T_46) begin
      wr_addr_reg_bits_1 <= _T_45;
    end
    if (reset) begin
      wr_addr_reg_bits_0 <= 16'h0;
    end else if (_T_43) begin
      wr_addr_reg_bits_0 <= 16'h0;
    end else if (_T_41) begin
      wr_addr_reg_bits_0 <= _T_40;
    end
    if (reset) begin
      wr_data_reg_valid <= 1'h0;
    end else begin
      wr_data_reg_valid <= io_wr_data_valid;
    end
    if (reset) begin
      wr_data_reg_bits <= 128'h0;
    end else begin
      wr_data_reg_bits <= io_wr_data_bits;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_63) begin
          $fwrite(32'h80000002,"wr_addr:%d %d, wr_data: %d, rd_addr:%d %d, rd_data: %d %d\n",mem_wr_addr,wr_addr_reg_valid,wr_data_reg_bits,mem_rd_addr,rd_addr_reg_valid,io_rd_data_valid,io_rd_data_bits); // @[mem.scala 167:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module MultiDimTime_105(
  input        clock,
  input        reset,
  input        io_in,
  output [1:0] io_out_0,
  output [1:0] io_out_1,
  output [1:0] io_out_2
);
  reg [15:0] regs_0; // @[mem.scala 67:12]
  reg [31:0] _RAND_0;
  reg [15:0] regs_1; // @[mem.scala 67:12]
  reg [31:0] _RAND_1;
  reg [15:0] regs_2; // @[mem.scala 67:12]
  reg [31:0] _RAND_2;
  wire [15:0] _GEN_10 = {{15'd0}, io_in}; // @[mem.scala 69:42]
  wire [15:0] _T_1 = regs_0 + _GEN_10; // @[mem.scala 69:42]
  wire  back_0 = _T_1 == 16'hc; // @[mem.scala 69:48]
  wire [15:0] _T_3 = regs_1 + _GEN_10; // @[mem.scala 69:42]
  wire  next_1 = _T_3 == 16'h16; // @[mem.scala 69:48]
  wire [15:0] _T_5 = regs_2 + _GEN_10; // @[mem.scala 69:42]
  wire  next_2 = _T_5 == 16'h10; // @[mem.scala 69:48]
  wire  back_1 = back_0 & next_1; // @[mem.scala 71:32]
  wire  back_2 = back_1 & next_2; // @[mem.scala 71:32]
  wire  _GEN_1 = back_0 ? 1'h0 : io_in; // @[mem.scala 90:20]
  wire  _GEN_3 = back_1 ? 1'h0 : 1'h1; // @[mem.scala 79:22]
  wire  _GEN_7 = back_2 ? 1'h0 : 1'h1; // @[mem.scala 79:22]
  assign io_out_0 = {{1'd0}, _GEN_1}; // @[mem.scala 92:19 mem.scala 95:19]
  assign io_out_1 = back_0 ? {{1'd0}, _GEN_3} : 2'h2; // @[mem.scala 81:21 mem.scala 84:21 mem.scala 87:19]
  assign io_out_2 = back_1 ? {{1'd0}, _GEN_7} : 2'h2; // @[mem.scala 81:21 mem.scala 84:21 mem.scala 87:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 16'h0;
    end else if (back_0) begin
      regs_0 <= 16'h0;
    end else begin
      regs_0 <= _T_1;
    end
    if (reset) begin
      regs_1 <= 16'h0;
    end else if (back_0) begin
      if (back_1) begin
        regs_1 <= 16'h0;
      end else begin
        regs_1 <= _T_3;
      end
    end
    if (reset) begin
      regs_2 <= 16'h0;
    end else if (back_1) begin
      if (back_2) begin
        regs_2 <= 16'h0;
      end else begin
        regs_2 <= _T_5;
      end
    end
  end
endmodule
module MemController_52(
  input          clock,
  input          reset,
  input          io_rd_valid,
  input          io_wr_valid,
  output         io_rd_data_valid,
  output [127:0] io_rd_data_bits,
  input          io_wr_data_valid,
  input  [127:0] io_wr_data_bits
);
  wire  MultiDimMem_clock; // @[mem.scala 31:19]
  wire  MultiDimMem_reset; // @[mem.scala 31:19]
  wire  MultiDimMem_io_rd_addr_valid; // @[mem.scala 31:19]
  wire [1:0] MultiDimMem_io_rd_addr_bits_0; // @[mem.scala 31:19]
  wire [1:0] MultiDimMem_io_rd_addr_bits_1; // @[mem.scala 31:19]
  wire [1:0] MultiDimMem_io_rd_addr_bits_2; // @[mem.scala 31:19]
  wire  MultiDimMem_io_rd_data_valid; // @[mem.scala 31:19]
  wire [127:0] MultiDimMem_io_rd_data_bits; // @[mem.scala 31:19]
  wire  MultiDimMem_io_wr_addr_valid; // @[mem.scala 31:19]
  wire [1:0] MultiDimMem_io_wr_addr_bits_0; // @[mem.scala 31:19]
  wire [1:0] MultiDimMem_io_wr_addr_bits_1; // @[mem.scala 31:19]
  wire [1:0] MultiDimMem_io_wr_addr_bits_2; // @[mem.scala 31:19]
  wire  MultiDimMem_io_wr_data_valid; // @[mem.scala 31:19]
  wire [127:0] MultiDimMem_io_wr_data_bits; // @[mem.scala 31:19]
  wire  MultiDimTime_clock; // @[mem.scala 32:23]
  wire  MultiDimTime_reset; // @[mem.scala 32:23]
  wire  MultiDimTime_io_in; // @[mem.scala 32:23]
  wire [1:0] MultiDimTime_io_out_0; // @[mem.scala 32:23]
  wire [1:0] MultiDimTime_io_out_1; // @[mem.scala 32:23]
  wire [1:0] MultiDimTime_io_out_2; // @[mem.scala 32:23]
  wire  MultiDimTime_1_clock; // @[mem.scala 33:23]
  wire  MultiDimTime_1_reset; // @[mem.scala 33:23]
  wire  MultiDimTime_1_io_in; // @[mem.scala 33:23]
  wire [1:0] MultiDimTime_1_io_out_0; // @[mem.scala 33:23]
  wire [1:0] MultiDimTime_1_io_out_1; // @[mem.scala 33:23]
  wire [1:0] MultiDimTime_1_io_out_2; // @[mem.scala 33:23]
  MultiDimMem_52 MultiDimMem ( // @[mem.scala 31:19]
    .clock(MultiDimMem_clock),
    .reset(MultiDimMem_reset),
    .io_rd_addr_valid(MultiDimMem_io_rd_addr_valid),
    .io_rd_addr_bits_0(MultiDimMem_io_rd_addr_bits_0),
    .io_rd_addr_bits_1(MultiDimMem_io_rd_addr_bits_1),
    .io_rd_addr_bits_2(MultiDimMem_io_rd_addr_bits_2),
    .io_rd_data_valid(MultiDimMem_io_rd_data_valid),
    .io_rd_data_bits(MultiDimMem_io_rd_data_bits),
    .io_wr_addr_valid(MultiDimMem_io_wr_addr_valid),
    .io_wr_addr_bits_0(MultiDimMem_io_wr_addr_bits_0),
    .io_wr_addr_bits_1(MultiDimMem_io_wr_addr_bits_1),
    .io_wr_addr_bits_2(MultiDimMem_io_wr_addr_bits_2),
    .io_wr_data_valid(MultiDimMem_io_wr_data_valid),
    .io_wr_data_bits(MultiDimMem_io_wr_data_bits)
  );
  MultiDimTime_105 MultiDimTime ( // @[mem.scala 32:23]
    .clock(MultiDimTime_clock),
    .reset(MultiDimTime_reset),
    .io_in(MultiDimTime_io_in),
    .io_out_0(MultiDimTime_io_out_0),
    .io_out_1(MultiDimTime_io_out_1),
    .io_out_2(MultiDimTime_io_out_2)
  );
  MultiDimTime_105 MultiDimTime_1 ( // @[mem.scala 33:23]
    .clock(MultiDimTime_1_clock),
    .reset(MultiDimTime_1_reset),
    .io_in(MultiDimTime_1_io_in),
    .io_out_0(MultiDimTime_1_io_out_0),
    .io_out_1(MultiDimTime_1_io_out_1),
    .io_out_2(MultiDimTime_1_io_out_2)
  );
  assign io_rd_data_valid = MultiDimMem_io_rd_data_valid; // @[mem.scala 50:14]
  assign io_rd_data_bits = MultiDimMem_io_rd_data_bits; // @[mem.scala 50:14]
  assign MultiDimMem_clock = clock;
  assign MultiDimMem_reset = reset;
  assign MultiDimMem_io_rd_addr_valid = io_rd_valid; // @[mem.scala 47:21]
  assign MultiDimMem_io_rd_addr_bits_0 = MultiDimTime_1_io_out_0; // @[mem.scala 46:20]
  assign MultiDimMem_io_rd_addr_bits_1 = MultiDimTime_1_io_out_1; // @[mem.scala 46:20]
  assign MultiDimMem_io_rd_addr_bits_2 = MultiDimTime_1_io_out_2; // @[mem.scala 46:20]
  assign MultiDimMem_io_wr_addr_valid = io_wr_valid; // @[mem.scala 43:21]
  assign MultiDimMem_io_wr_addr_bits_0 = MultiDimTime_io_out_0; // @[mem.scala 42:20]
  assign MultiDimMem_io_wr_addr_bits_1 = MultiDimTime_io_out_1; // @[mem.scala 42:20]
  assign MultiDimMem_io_wr_addr_bits_2 = MultiDimTime_io_out_2; // @[mem.scala 42:20]
  assign MultiDimMem_io_wr_data_valid = io_wr_data_valid; // @[mem.scala 51:15]
  assign MultiDimMem_io_wr_data_bits = io_wr_data_bits; // @[mem.scala 51:15]
  assign MultiDimTime_clock = clock;
  assign MultiDimTime_reset = reset;
  assign MultiDimTime_io_in = io_wr_valid; // @[mem.scala 41:14]
  assign MultiDimTime_1_clock = clock;
  assign MultiDimTime_1_reset = reset;
  assign MultiDimTime_1_io_in = io_rd_valid; // @[mem.scala 45:14]
endmodule
module PEArray2D(
  input          clock,
  input          reset,
  output         io_data_2_out_0_valid,
  output [127:0] io_data_2_out_0_bits,
  output         io_data_2_out_1_valid,
  output [127:0] io_data_2_out_1_bits,
  output         io_data_2_out_2_valid,
  output [127:0] io_data_2_out_2_bits,
  output         io_data_2_out_3_valid,
  output [127:0] io_data_2_out_3_bits,
  output         io_data_2_out_4_valid,
  output [127:0] io_data_2_out_4_bits,
  output         io_data_2_out_5_valid,
  output [127:0] io_data_2_out_5_bits,
  output         io_data_2_out_6_valid,
  output [127:0] io_data_2_out_6_bits,
  output         io_data_2_out_7_valid,
  output [127:0] io_data_2_out_7_bits,
  output         io_data_2_out_8_valid,
  output [127:0] io_data_2_out_8_bits,
  output         io_data_2_out_9_valid,
  output [127:0] io_data_2_out_9_bits,
  output         io_data_2_out_10_valid,
  output [127:0] io_data_2_out_10_bits,
  output         io_data_2_out_11_valid,
  output [127:0] io_data_2_out_11_bits,
  output         io_data_2_out_12_valid,
  output [127:0] io_data_2_out_12_bits,
  output         io_data_2_out_13_valid,
  output [127:0] io_data_2_out_13_bits,
  output         io_data_2_out_14_valid,
  output [127:0] io_data_2_out_14_bits,
  output         io_data_2_out_15_valid,
  output [127:0] io_data_2_out_15_bits,
  output         io_data_2_out_16_valid,
  output [127:0] io_data_2_out_16_bits,
  output         io_data_2_out_17_valid,
  output [127:0] io_data_2_out_17_bits,
  output         io_data_2_out_18_valid,
  output [127:0] io_data_2_out_18_bits,
  output         io_data_2_out_19_valid,
  output [127:0] io_data_2_out_19_bits,
  output         io_data_2_out_20_valid,
  output [127:0] io_data_2_out_20_bits,
  output         io_data_2_out_21_valid,
  output [127:0] io_data_2_out_21_bits,
  output         io_data_2_out_22_valid,
  output [127:0] io_data_2_out_22_bits,
  output         io_data_2_out_23_valid,
  output [127:0] io_data_2_out_23_bits,
  output         io_data_2_out_24_valid,
  output [127:0] io_data_2_out_24_bits,
  output         io_data_2_out_25_valid,
  output [127:0] io_data_2_out_25_bits,
  output         io_data_2_out_26_valid,
  output [127:0] io_data_2_out_26_bits,
  output         io_data_2_out_27_valid,
  output [127:0] io_data_2_out_27_bits,
  output         io_data_2_out_28_valid,
  output [127:0] io_data_2_out_28_bits,
  output         io_data_2_out_29_valid,
  output [127:0] io_data_2_out_29_bits,
  input          io_data_1_in_0_valid,
  input          io_data_1_in_0_bits_valid,
  input  [127:0] io_data_1_in_0_bits_bits,
  input          io_data_1_in_1_valid,
  input          io_data_1_in_1_bits_valid,
  input  [127:0] io_data_1_in_1_bits_bits,
  input          io_data_1_in_2_valid,
  input          io_data_1_in_2_bits_valid,
  input  [127:0] io_data_1_in_2_bits_bits,
  input          io_data_1_in_3_valid,
  input          io_data_1_in_3_bits_valid,
  input  [127:0] io_data_1_in_3_bits_bits,
  input          io_data_1_in_4_valid,
  input          io_data_1_in_4_bits_valid,
  input  [127:0] io_data_1_in_4_bits_bits,
  input          io_data_1_in_5_valid,
  input          io_data_1_in_5_bits_valid,
  input  [127:0] io_data_1_in_5_bits_bits,
  input          io_data_1_in_6_valid,
  input          io_data_1_in_6_bits_valid,
  input  [127:0] io_data_1_in_6_bits_bits,
  input          io_data_1_in_7_valid,
  input          io_data_1_in_7_bits_valid,
  input  [127:0] io_data_1_in_7_bits_bits,
  input          io_data_1_in_8_valid,
  input          io_data_1_in_8_bits_valid,
  input  [127:0] io_data_1_in_8_bits_bits,
  input          io_data_1_in_9_valid,
  input          io_data_1_in_9_bits_valid,
  input  [127:0] io_data_1_in_9_bits_bits,
  input          io_data_1_in_10_valid,
  input          io_data_1_in_10_bits_valid,
  input  [127:0] io_data_1_in_10_bits_bits,
  input          io_data_1_in_11_valid,
  input          io_data_1_in_11_bits_valid,
  input  [127:0] io_data_1_in_11_bits_bits,
  input          io_data_1_in_12_valid,
  input          io_data_1_in_12_bits_valid,
  input  [127:0] io_data_1_in_12_bits_bits,
  input          io_data_1_in_13_valid,
  input          io_data_1_in_13_bits_valid,
  input  [127:0] io_data_1_in_13_bits_bits,
  input          io_data_1_in_14_valid,
  input          io_data_1_in_14_bits_valid,
  input  [127:0] io_data_1_in_14_bits_bits,
  input          io_data_1_in_15_valid,
  input          io_data_1_in_15_bits_valid,
  input  [127:0] io_data_1_in_15_bits_bits,
  input          io_data_1_in_16_valid,
  input          io_data_1_in_16_bits_valid,
  input  [127:0] io_data_1_in_16_bits_bits,
  input          io_data_1_in_17_valid,
  input          io_data_1_in_17_bits_valid,
  input  [127:0] io_data_1_in_17_bits_bits,
  input          io_data_1_in_18_valid,
  input          io_data_1_in_18_bits_valid,
  input  [127:0] io_data_1_in_18_bits_bits,
  input          io_data_1_in_19_valid,
  input          io_data_1_in_19_bits_valid,
  input  [127:0] io_data_1_in_19_bits_bits,
  input          io_data_1_in_20_valid,
  input          io_data_1_in_20_bits_valid,
  input  [127:0] io_data_1_in_20_bits_bits,
  input          io_data_1_in_21_valid,
  input          io_data_1_in_21_bits_valid,
  input  [127:0] io_data_1_in_21_bits_bits,
  input          io_data_1_in_22_valid,
  input          io_data_1_in_22_bits_valid,
  input  [127:0] io_data_1_in_22_bits_bits,
  input          io_data_1_in_23_valid,
  input          io_data_1_in_23_bits_valid,
  input  [127:0] io_data_1_in_23_bits_bits,
  input          io_data_1_in_24_valid,
  input          io_data_1_in_24_bits_valid,
  input  [127:0] io_data_1_in_24_bits_bits,
  input          io_data_1_in_25_valid,
  input          io_data_1_in_25_bits_valid,
  input  [127:0] io_data_1_in_25_bits_bits,
  input          io_data_1_in_26_valid,
  input          io_data_1_in_26_bits_valid,
  input  [127:0] io_data_1_in_26_bits_bits,
  input          io_data_1_in_27_valid,
  input          io_data_1_in_27_bits_valid,
  input  [127:0] io_data_1_in_27_bits_bits,
  input          io_data_1_in_28_valid,
  input          io_data_1_in_28_bits_valid,
  input  [127:0] io_data_1_in_28_bits_bits,
  input          io_data_1_in_29_valid,
  input          io_data_1_in_29_bits_valid,
  input  [127:0] io_data_1_in_29_bits_bits,
  input          io_data_0_in_0_valid,
  input          io_data_0_in_0_bits_valid,
  input  [15:0]  io_data_0_in_0_bits_bits,
  input          io_data_0_in_1_valid,
  input          io_data_0_in_1_bits_valid,
  input  [15:0]  io_data_0_in_1_bits_bits,
  input          io_data_0_in_2_valid,
  input          io_data_0_in_2_bits_valid,
  input  [15:0]  io_data_0_in_2_bits_bits,
  input          io_data_0_in_3_valid,
  input          io_data_0_in_3_bits_valid,
  input  [15:0]  io_data_0_in_3_bits_bits,
  input          io_data_0_in_4_valid,
  input          io_data_0_in_4_bits_valid,
  input  [15:0]  io_data_0_in_4_bits_bits,
  input          io_data_0_in_5_valid,
  input          io_data_0_in_5_bits_valid,
  input  [15:0]  io_data_0_in_5_bits_bits,
  input          io_data_0_in_6_valid,
  input          io_data_0_in_6_bits_valid,
  input  [15:0]  io_data_0_in_6_bits_bits,
  input          io_data_0_in_7_valid,
  input          io_data_0_in_7_bits_valid,
  input  [15:0]  io_data_0_in_7_bits_bits,
  input          io_data_0_in_8_valid,
  input          io_data_0_in_8_bits_valid,
  input  [15:0]  io_data_0_in_8_bits_bits,
  input          io_data_0_in_9_valid,
  input          io_data_0_in_9_bits_valid,
  input  [15:0]  io_data_0_in_9_bits_bits,
  input          io_data_0_in_10_valid,
  input          io_data_0_in_10_bits_valid,
  input  [15:0]  io_data_0_in_10_bits_bits,
  input          io_data_0_in_11_valid,
  input          io_data_0_in_11_bits_valid,
  input  [15:0]  io_data_0_in_11_bits_bits,
  input          io_data_0_in_12_valid,
  input          io_data_0_in_12_bits_valid,
  input  [15:0]  io_data_0_in_12_bits_bits,
  input          io_data_0_in_13_valid,
  input          io_data_0_in_13_bits_valid,
  input  [15:0]  io_data_0_in_13_bits_bits,
  input          io_data_0_in_14_valid,
  input          io_data_0_in_14_bits_valid,
  input  [15:0]  io_data_0_in_14_bits_bits,
  input          io_data_0_in_15_valid,
  input          io_data_0_in_15_bits_valid,
  input  [15:0]  io_data_0_in_15_bits_bits,
  input          io_data_0_in_16_valid,
  input          io_data_0_in_16_bits_valid,
  input  [15:0]  io_data_0_in_16_bits_bits,
  input          io_data_0_in_17_valid,
  input          io_data_0_in_17_bits_valid,
  input  [15:0]  io_data_0_in_17_bits_bits,
  input          io_data_0_in_18_valid,
  input          io_data_0_in_18_bits_valid,
  input  [15:0]  io_data_0_in_18_bits_bits,
  input          io_data_0_in_19_valid,
  input          io_data_0_in_19_bits_valid,
  input  [15:0]  io_data_0_in_19_bits_bits,
  input          io_data_0_in_20_valid,
  input          io_data_0_in_20_bits_valid,
  input  [15:0]  io_data_0_in_20_bits_bits,
  input          io_data_0_in_21_valid,
  input          io_data_0_in_21_bits_valid,
  input  [15:0]  io_data_0_in_21_bits_bits,
  input          io_exec_valid,
  input          io_out_valid
);
  wire  MultiDimTime_clock; // @[pe.scala 165:25]
  wire  MultiDimTime_reset; // @[pe.scala 165:25]
  wire  MultiDimTime_io_in; // @[pe.scala 165:25]
  wire [1:0] MultiDimTime_io_out_0; // @[pe.scala 165:25]
  wire [1:0] MultiDimTime_io_out_1; // @[pe.scala 165:25]
  wire [1:0] MultiDimTime_io_out_2; // @[pe.scala 165:25]
  wire [15:0] MultiDimTime_io_index_0; // @[pe.scala 165:25]
  wire [15:0] MultiDimTime_io_index_1; // @[pe.scala 165:25]
  wire [15:0] MultiDimTime_io_index_2; // @[pe.scala 165:25]
  wire  PE_clock; // @[pe.scala 187:13]
  wire  PE_reset; // @[pe.scala 187:13]
  wire  PE_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_1_clock; // @[pe.scala 187:13]
  wire  PE_1_reset; // @[pe.scala 187:13]
  wire  PE_1_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_1_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_1_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_1_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_1_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_1_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_1_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_1_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_1_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_1_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_1_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_2_clock; // @[pe.scala 187:13]
  wire  PE_2_reset; // @[pe.scala 187:13]
  wire  PE_2_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_2_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_2_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_2_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_2_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_2_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_2_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_2_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_2_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_2_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_2_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_3_clock; // @[pe.scala 187:13]
  wire  PE_3_reset; // @[pe.scala 187:13]
  wire  PE_3_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_3_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_3_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_3_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_3_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_3_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_3_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_3_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_3_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_3_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_3_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_4_clock; // @[pe.scala 187:13]
  wire  PE_4_reset; // @[pe.scala 187:13]
  wire  PE_4_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_4_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_4_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_4_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_4_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_4_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_4_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_4_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_4_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_4_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_4_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_5_clock; // @[pe.scala 187:13]
  wire  PE_5_reset; // @[pe.scala 187:13]
  wire  PE_5_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_5_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_5_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_5_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_5_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_5_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_5_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_5_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_5_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_5_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_5_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_6_clock; // @[pe.scala 187:13]
  wire  PE_6_reset; // @[pe.scala 187:13]
  wire  PE_6_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_6_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_6_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_6_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_6_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_6_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_6_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_6_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_6_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_6_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_6_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_7_clock; // @[pe.scala 187:13]
  wire  PE_7_reset; // @[pe.scala 187:13]
  wire  PE_7_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_7_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_7_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_7_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_7_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_7_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_7_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_7_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_7_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_7_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_7_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_8_clock; // @[pe.scala 187:13]
  wire  PE_8_reset; // @[pe.scala 187:13]
  wire  PE_8_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_8_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_8_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_8_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_8_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_8_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_8_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_8_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_8_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_8_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_8_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_9_clock; // @[pe.scala 187:13]
  wire  PE_9_reset; // @[pe.scala 187:13]
  wire  PE_9_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_9_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_9_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_9_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_9_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_9_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_9_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_9_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_9_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_9_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_9_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_10_clock; // @[pe.scala 187:13]
  wire  PE_10_reset; // @[pe.scala 187:13]
  wire  PE_10_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_10_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_10_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_10_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_10_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_10_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_10_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_10_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_10_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_10_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_10_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_11_clock; // @[pe.scala 187:13]
  wire  PE_11_reset; // @[pe.scala 187:13]
  wire  PE_11_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_11_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_11_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_11_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_11_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_11_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_11_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_11_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_11_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_11_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_11_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_12_clock; // @[pe.scala 187:13]
  wire  PE_12_reset; // @[pe.scala 187:13]
  wire  PE_12_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_12_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_12_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_12_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_12_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_12_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_12_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_12_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_12_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_12_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_12_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_13_clock; // @[pe.scala 187:13]
  wire  PE_13_reset; // @[pe.scala 187:13]
  wire  PE_13_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_13_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_13_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_13_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_13_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_13_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_13_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_13_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_13_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_13_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_13_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_14_clock; // @[pe.scala 187:13]
  wire  PE_14_reset; // @[pe.scala 187:13]
  wire  PE_14_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_14_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_14_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_14_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_14_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_14_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_14_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_14_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_14_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_14_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_14_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_15_clock; // @[pe.scala 187:13]
  wire  PE_15_reset; // @[pe.scala 187:13]
  wire  PE_15_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_15_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_15_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_15_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_15_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_15_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_15_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_15_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_15_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_15_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_15_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_16_clock; // @[pe.scala 187:13]
  wire  PE_16_reset; // @[pe.scala 187:13]
  wire  PE_16_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_16_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_16_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_16_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_16_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_16_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_16_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_16_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_16_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_16_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_16_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_17_clock; // @[pe.scala 187:13]
  wire  PE_17_reset; // @[pe.scala 187:13]
  wire  PE_17_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_17_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_17_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_17_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_17_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_17_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_17_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_17_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_17_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_17_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_17_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_18_clock; // @[pe.scala 187:13]
  wire  PE_18_reset; // @[pe.scala 187:13]
  wire  PE_18_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_18_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_18_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_18_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_18_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_18_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_18_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_18_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_18_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_18_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_18_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_19_clock; // @[pe.scala 187:13]
  wire  PE_19_reset; // @[pe.scala 187:13]
  wire  PE_19_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_19_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_19_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_19_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_19_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_19_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_19_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_19_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_19_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_19_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_19_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_20_clock; // @[pe.scala 187:13]
  wire  PE_20_reset; // @[pe.scala 187:13]
  wire  PE_20_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_20_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_20_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_20_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_20_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_20_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_20_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_20_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_20_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_20_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_20_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_21_clock; // @[pe.scala 187:13]
  wire  PE_21_reset; // @[pe.scala 187:13]
  wire  PE_21_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_21_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_21_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_21_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_21_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_21_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_21_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_21_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_21_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_21_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_21_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_22_clock; // @[pe.scala 187:13]
  wire  PE_22_reset; // @[pe.scala 187:13]
  wire  PE_22_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_22_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_22_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_22_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_22_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_22_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_22_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_22_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_22_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_22_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_22_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_23_clock; // @[pe.scala 187:13]
  wire  PE_23_reset; // @[pe.scala 187:13]
  wire  PE_23_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_23_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_23_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_23_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_23_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_23_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_23_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_23_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_23_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_23_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_23_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_24_clock; // @[pe.scala 187:13]
  wire  PE_24_reset; // @[pe.scala 187:13]
  wire  PE_24_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_24_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_24_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_24_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_24_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_24_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_24_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_24_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_24_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_24_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_24_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_25_clock; // @[pe.scala 187:13]
  wire  PE_25_reset; // @[pe.scala 187:13]
  wire  PE_25_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_25_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_25_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_25_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_25_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_25_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_25_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_25_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_25_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_25_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_25_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_26_clock; // @[pe.scala 187:13]
  wire  PE_26_reset; // @[pe.scala 187:13]
  wire  PE_26_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_26_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_26_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_26_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_26_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_26_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_26_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_26_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_26_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_26_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_26_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_27_clock; // @[pe.scala 187:13]
  wire  PE_27_reset; // @[pe.scala 187:13]
  wire  PE_27_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_27_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_27_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_27_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_27_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_27_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_27_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_27_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_27_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_27_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_27_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_28_clock; // @[pe.scala 187:13]
  wire  PE_28_reset; // @[pe.scala 187:13]
  wire  PE_28_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_28_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_28_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_28_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_28_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_28_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_28_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_28_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_28_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_28_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_28_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_29_clock; // @[pe.scala 187:13]
  wire  PE_29_reset; // @[pe.scala 187:13]
  wire  PE_29_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_29_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_29_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_29_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_29_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_29_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_29_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_29_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_29_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_29_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_29_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_30_clock; // @[pe.scala 187:13]
  wire  PE_30_reset; // @[pe.scala 187:13]
  wire  PE_30_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_30_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_30_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_30_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_30_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_30_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_30_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_30_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_30_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_30_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_30_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_31_clock; // @[pe.scala 187:13]
  wire  PE_31_reset; // @[pe.scala 187:13]
  wire  PE_31_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_31_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_31_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_31_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_31_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_31_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_31_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_31_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_31_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_31_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_31_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_32_clock; // @[pe.scala 187:13]
  wire  PE_32_reset; // @[pe.scala 187:13]
  wire  PE_32_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_32_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_32_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_32_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_32_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_32_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_32_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_32_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_32_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_32_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_32_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_33_clock; // @[pe.scala 187:13]
  wire  PE_33_reset; // @[pe.scala 187:13]
  wire  PE_33_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_33_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_33_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_33_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_33_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_33_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_33_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_33_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_33_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_33_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_33_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_34_clock; // @[pe.scala 187:13]
  wire  PE_34_reset; // @[pe.scala 187:13]
  wire  PE_34_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_34_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_34_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_34_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_34_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_34_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_34_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_34_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_34_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_34_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_34_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_35_clock; // @[pe.scala 187:13]
  wire  PE_35_reset; // @[pe.scala 187:13]
  wire  PE_35_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_35_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_35_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_35_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_35_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_35_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_35_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_35_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_35_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_35_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_35_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_36_clock; // @[pe.scala 187:13]
  wire  PE_36_reset; // @[pe.scala 187:13]
  wire  PE_36_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_36_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_36_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_36_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_36_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_36_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_36_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_36_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_36_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_36_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_36_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_37_clock; // @[pe.scala 187:13]
  wire  PE_37_reset; // @[pe.scala 187:13]
  wire  PE_37_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_37_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_37_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_37_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_37_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_37_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_37_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_37_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_37_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_37_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_37_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_38_clock; // @[pe.scala 187:13]
  wire  PE_38_reset; // @[pe.scala 187:13]
  wire  PE_38_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_38_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_38_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_38_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_38_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_38_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_38_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_38_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_38_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_38_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_38_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_39_clock; // @[pe.scala 187:13]
  wire  PE_39_reset; // @[pe.scala 187:13]
  wire  PE_39_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_39_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_39_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_39_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_39_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_39_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_39_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_39_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_39_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_39_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_39_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_40_clock; // @[pe.scala 187:13]
  wire  PE_40_reset; // @[pe.scala 187:13]
  wire  PE_40_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_40_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_40_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_40_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_40_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_40_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_40_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_40_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_40_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_40_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_40_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_41_clock; // @[pe.scala 187:13]
  wire  PE_41_reset; // @[pe.scala 187:13]
  wire  PE_41_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_41_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_41_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_41_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_41_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_41_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_41_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_41_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_41_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_41_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_41_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_42_clock; // @[pe.scala 187:13]
  wire  PE_42_reset; // @[pe.scala 187:13]
  wire  PE_42_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_42_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_42_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_42_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_42_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_42_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_42_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_42_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_42_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_42_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_42_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_43_clock; // @[pe.scala 187:13]
  wire  PE_43_reset; // @[pe.scala 187:13]
  wire  PE_43_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_43_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_43_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_43_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_43_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_43_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_43_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_43_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_43_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_43_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_43_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_44_clock; // @[pe.scala 187:13]
  wire  PE_44_reset; // @[pe.scala 187:13]
  wire  PE_44_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_44_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_44_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_44_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_44_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_44_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_44_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_44_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_44_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_44_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_44_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_45_clock; // @[pe.scala 187:13]
  wire  PE_45_reset; // @[pe.scala 187:13]
  wire  PE_45_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_45_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_45_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_45_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_45_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_45_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_45_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_45_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_45_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_45_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_45_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_46_clock; // @[pe.scala 187:13]
  wire  PE_46_reset; // @[pe.scala 187:13]
  wire  PE_46_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_46_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_46_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_46_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_46_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_46_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_46_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_46_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_46_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_46_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_46_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_47_clock; // @[pe.scala 187:13]
  wire  PE_47_reset; // @[pe.scala 187:13]
  wire  PE_47_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_47_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_47_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_47_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_47_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_47_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_47_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_47_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_47_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_47_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_47_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_48_clock; // @[pe.scala 187:13]
  wire  PE_48_reset; // @[pe.scala 187:13]
  wire  PE_48_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_48_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_48_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_48_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_48_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_48_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_48_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_48_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_48_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_48_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_48_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_49_clock; // @[pe.scala 187:13]
  wire  PE_49_reset; // @[pe.scala 187:13]
  wire  PE_49_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_49_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_49_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_49_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_49_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_49_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_49_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_49_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_49_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_49_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_49_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_50_clock; // @[pe.scala 187:13]
  wire  PE_50_reset; // @[pe.scala 187:13]
  wire  PE_50_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_50_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_50_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_50_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_50_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_50_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_50_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_50_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_50_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_50_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_50_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_51_clock; // @[pe.scala 187:13]
  wire  PE_51_reset; // @[pe.scala 187:13]
  wire  PE_51_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_51_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_51_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_51_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_51_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_51_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_51_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_51_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_51_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_51_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_51_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_52_clock; // @[pe.scala 187:13]
  wire  PE_52_reset; // @[pe.scala 187:13]
  wire  PE_52_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_52_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_52_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_52_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_52_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_52_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_52_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_52_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_52_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_52_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_52_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_53_clock; // @[pe.scala 187:13]
  wire  PE_53_reset; // @[pe.scala 187:13]
  wire  PE_53_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_53_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_53_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_53_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_53_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_53_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_53_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_53_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_53_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_53_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_53_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_54_clock; // @[pe.scala 187:13]
  wire  PE_54_reset; // @[pe.scala 187:13]
  wire  PE_54_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_54_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_54_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_54_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_54_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_54_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_54_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_54_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_54_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_54_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_54_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_55_clock; // @[pe.scala 187:13]
  wire  PE_55_reset; // @[pe.scala 187:13]
  wire  PE_55_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_55_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_55_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_55_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_55_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_55_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_55_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_55_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_55_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_55_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_55_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_56_clock; // @[pe.scala 187:13]
  wire  PE_56_reset; // @[pe.scala 187:13]
  wire  PE_56_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_56_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_56_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_56_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_56_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_56_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_56_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_56_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_56_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_56_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_56_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_57_clock; // @[pe.scala 187:13]
  wire  PE_57_reset; // @[pe.scala 187:13]
  wire  PE_57_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_57_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_57_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_57_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_57_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_57_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_57_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_57_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_57_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_57_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_57_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_58_clock; // @[pe.scala 187:13]
  wire  PE_58_reset; // @[pe.scala 187:13]
  wire  PE_58_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_58_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_58_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_58_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_58_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_58_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_58_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_58_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_58_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_58_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_58_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_59_clock; // @[pe.scala 187:13]
  wire  PE_59_reset; // @[pe.scala 187:13]
  wire  PE_59_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_59_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_59_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_59_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_59_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_59_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_59_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_59_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_59_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_59_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_59_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_60_clock; // @[pe.scala 187:13]
  wire  PE_60_reset; // @[pe.scala 187:13]
  wire  PE_60_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_60_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_60_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_60_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_60_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_60_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_60_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_60_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_60_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_60_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_60_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_61_clock; // @[pe.scala 187:13]
  wire  PE_61_reset; // @[pe.scala 187:13]
  wire  PE_61_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_61_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_61_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_61_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_61_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_61_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_61_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_61_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_61_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_61_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_61_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_62_clock; // @[pe.scala 187:13]
  wire  PE_62_reset; // @[pe.scala 187:13]
  wire  PE_62_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_62_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_62_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_62_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_62_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_62_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_62_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_62_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_62_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_62_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_62_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_63_clock; // @[pe.scala 187:13]
  wire  PE_63_reset; // @[pe.scala 187:13]
  wire  PE_63_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_63_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_63_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_63_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_63_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_63_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_63_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_63_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_63_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_63_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_63_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_64_clock; // @[pe.scala 187:13]
  wire  PE_64_reset; // @[pe.scala 187:13]
  wire  PE_64_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_64_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_64_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_64_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_64_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_64_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_64_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_64_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_64_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_64_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_64_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_65_clock; // @[pe.scala 187:13]
  wire  PE_65_reset; // @[pe.scala 187:13]
  wire  PE_65_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_65_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_65_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_65_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_65_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_65_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_65_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_65_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_65_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_65_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_65_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_66_clock; // @[pe.scala 187:13]
  wire  PE_66_reset; // @[pe.scala 187:13]
  wire  PE_66_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_66_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_66_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_66_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_66_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_66_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_66_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_66_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_66_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_66_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_66_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_67_clock; // @[pe.scala 187:13]
  wire  PE_67_reset; // @[pe.scala 187:13]
  wire  PE_67_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_67_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_67_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_67_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_67_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_67_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_67_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_67_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_67_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_67_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_67_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_68_clock; // @[pe.scala 187:13]
  wire  PE_68_reset; // @[pe.scala 187:13]
  wire  PE_68_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_68_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_68_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_68_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_68_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_68_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_68_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_68_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_68_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_68_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_68_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_69_clock; // @[pe.scala 187:13]
  wire  PE_69_reset; // @[pe.scala 187:13]
  wire  PE_69_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_69_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_69_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_69_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_69_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_69_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_69_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_69_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_69_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_69_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_69_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_70_clock; // @[pe.scala 187:13]
  wire  PE_70_reset; // @[pe.scala 187:13]
  wire  PE_70_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_70_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_70_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_70_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_70_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_70_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_70_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_70_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_70_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_70_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_70_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_71_clock; // @[pe.scala 187:13]
  wire  PE_71_reset; // @[pe.scala 187:13]
  wire  PE_71_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_71_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_71_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_71_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_71_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_71_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_71_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_71_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_71_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_71_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_71_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_72_clock; // @[pe.scala 187:13]
  wire  PE_72_reset; // @[pe.scala 187:13]
  wire  PE_72_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_72_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_72_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_72_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_72_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_72_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_72_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_72_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_72_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_72_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_72_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_73_clock; // @[pe.scala 187:13]
  wire  PE_73_reset; // @[pe.scala 187:13]
  wire  PE_73_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_73_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_73_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_73_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_73_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_73_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_73_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_73_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_73_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_73_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_73_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_74_clock; // @[pe.scala 187:13]
  wire  PE_74_reset; // @[pe.scala 187:13]
  wire  PE_74_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_74_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_74_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_74_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_74_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_74_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_74_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_74_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_74_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_74_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_74_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_75_clock; // @[pe.scala 187:13]
  wire  PE_75_reset; // @[pe.scala 187:13]
  wire  PE_75_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_75_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_75_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_75_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_75_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_75_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_75_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_75_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_75_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_75_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_75_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_76_clock; // @[pe.scala 187:13]
  wire  PE_76_reset; // @[pe.scala 187:13]
  wire  PE_76_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_76_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_76_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_76_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_76_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_76_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_76_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_76_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_76_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_76_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_76_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_77_clock; // @[pe.scala 187:13]
  wire  PE_77_reset; // @[pe.scala 187:13]
  wire  PE_77_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_77_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_77_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_77_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_77_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_77_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_77_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_77_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_77_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_77_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_77_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_78_clock; // @[pe.scala 187:13]
  wire  PE_78_reset; // @[pe.scala 187:13]
  wire  PE_78_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_78_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_78_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_78_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_78_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_78_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_78_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_78_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_78_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_78_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_78_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_79_clock; // @[pe.scala 187:13]
  wire  PE_79_reset; // @[pe.scala 187:13]
  wire  PE_79_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_79_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_79_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_79_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_79_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_79_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_79_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_79_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_79_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_79_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_79_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_80_clock; // @[pe.scala 187:13]
  wire  PE_80_reset; // @[pe.scala 187:13]
  wire  PE_80_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_80_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_80_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_80_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_80_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_80_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_80_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_80_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_80_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_80_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_80_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_81_clock; // @[pe.scala 187:13]
  wire  PE_81_reset; // @[pe.scala 187:13]
  wire  PE_81_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_81_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_81_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_81_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_81_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_81_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_81_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_81_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_81_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_81_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_81_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_82_clock; // @[pe.scala 187:13]
  wire  PE_82_reset; // @[pe.scala 187:13]
  wire  PE_82_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_82_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_82_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_82_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_82_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_82_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_82_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_82_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_82_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_82_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_82_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_83_clock; // @[pe.scala 187:13]
  wire  PE_83_reset; // @[pe.scala 187:13]
  wire  PE_83_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_83_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_83_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_83_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_83_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_83_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_83_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_83_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_83_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_83_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_83_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_84_clock; // @[pe.scala 187:13]
  wire  PE_84_reset; // @[pe.scala 187:13]
  wire  PE_84_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_84_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_84_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_84_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_84_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_84_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_84_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_84_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_84_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_84_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_84_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_85_clock; // @[pe.scala 187:13]
  wire  PE_85_reset; // @[pe.scala 187:13]
  wire  PE_85_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_85_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_85_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_85_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_85_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_85_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_85_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_85_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_85_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_85_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_85_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_86_clock; // @[pe.scala 187:13]
  wire  PE_86_reset; // @[pe.scala 187:13]
  wire  PE_86_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_86_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_86_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_86_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_86_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_86_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_86_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_86_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_86_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_86_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_86_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_87_clock; // @[pe.scala 187:13]
  wire  PE_87_reset; // @[pe.scala 187:13]
  wire  PE_87_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_87_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_87_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_87_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_87_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_87_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_87_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_87_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_87_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_87_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_87_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_88_clock; // @[pe.scala 187:13]
  wire  PE_88_reset; // @[pe.scala 187:13]
  wire  PE_88_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_88_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_88_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_88_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_88_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_88_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_88_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_88_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_88_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_88_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_88_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_89_clock; // @[pe.scala 187:13]
  wire  PE_89_reset; // @[pe.scala 187:13]
  wire  PE_89_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_89_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_89_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_89_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_89_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_89_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_89_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_89_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_89_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_89_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_89_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_90_clock; // @[pe.scala 187:13]
  wire  PE_90_reset; // @[pe.scala 187:13]
  wire  PE_90_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_90_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_90_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_90_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_90_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_90_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_90_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_90_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_90_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_90_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_90_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_91_clock; // @[pe.scala 187:13]
  wire  PE_91_reset; // @[pe.scala 187:13]
  wire  PE_91_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_91_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_91_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_91_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_91_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_91_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_91_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_91_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_91_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_91_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_91_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_92_clock; // @[pe.scala 187:13]
  wire  PE_92_reset; // @[pe.scala 187:13]
  wire  PE_92_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_92_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_92_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_92_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_92_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_92_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_92_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_92_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_92_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_92_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_92_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_93_clock; // @[pe.scala 187:13]
  wire  PE_93_reset; // @[pe.scala 187:13]
  wire  PE_93_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_93_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_93_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_93_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_93_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_93_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_93_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_93_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_93_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_93_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_93_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_94_clock; // @[pe.scala 187:13]
  wire  PE_94_reset; // @[pe.scala 187:13]
  wire  PE_94_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_94_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_94_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_94_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_94_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_94_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_94_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_94_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_94_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_94_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_94_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_95_clock; // @[pe.scala 187:13]
  wire  PE_95_reset; // @[pe.scala 187:13]
  wire  PE_95_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_95_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_95_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_95_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_95_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_95_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_95_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_95_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_95_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_95_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_95_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_96_clock; // @[pe.scala 187:13]
  wire  PE_96_reset; // @[pe.scala 187:13]
  wire  PE_96_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_96_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_96_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_96_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_96_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_96_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_96_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_96_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_96_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_96_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_96_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_97_clock; // @[pe.scala 187:13]
  wire  PE_97_reset; // @[pe.scala 187:13]
  wire  PE_97_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_97_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_97_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_97_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_97_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_97_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_97_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_97_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_97_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_97_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_97_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_98_clock; // @[pe.scala 187:13]
  wire  PE_98_reset; // @[pe.scala 187:13]
  wire  PE_98_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_98_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_98_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_98_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_98_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_98_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_98_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_98_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_98_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_98_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_98_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_99_clock; // @[pe.scala 187:13]
  wire  PE_99_reset; // @[pe.scala 187:13]
  wire  PE_99_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_99_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_99_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_99_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_99_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_99_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_99_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_99_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_99_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_99_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_99_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_100_clock; // @[pe.scala 187:13]
  wire  PE_100_reset; // @[pe.scala 187:13]
  wire  PE_100_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_100_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_100_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_100_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_100_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_100_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_100_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_100_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_100_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_100_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_100_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_101_clock; // @[pe.scala 187:13]
  wire  PE_101_reset; // @[pe.scala 187:13]
  wire  PE_101_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_101_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_101_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_101_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_101_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_101_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_101_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_101_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_101_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_101_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_101_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_102_clock; // @[pe.scala 187:13]
  wire  PE_102_reset; // @[pe.scala 187:13]
  wire  PE_102_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_102_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_102_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_102_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_102_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_102_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_102_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_102_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_102_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_102_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_102_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_103_clock; // @[pe.scala 187:13]
  wire  PE_103_reset; // @[pe.scala 187:13]
  wire  PE_103_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_103_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_103_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_103_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_103_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_103_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_103_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_103_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_103_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_103_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_103_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_104_clock; // @[pe.scala 187:13]
  wire  PE_104_reset; // @[pe.scala 187:13]
  wire  PE_104_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_104_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_104_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_104_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_104_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_104_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_104_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_104_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_104_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_104_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_104_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_105_clock; // @[pe.scala 187:13]
  wire  PE_105_reset; // @[pe.scala 187:13]
  wire  PE_105_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_105_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_105_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_105_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_105_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_105_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_105_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_105_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_105_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_105_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_105_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_106_clock; // @[pe.scala 187:13]
  wire  PE_106_reset; // @[pe.scala 187:13]
  wire  PE_106_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_106_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_106_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_106_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_106_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_106_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_106_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_106_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_106_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_106_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_106_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_107_clock; // @[pe.scala 187:13]
  wire  PE_107_reset; // @[pe.scala 187:13]
  wire  PE_107_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_107_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_107_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_107_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_107_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_107_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_107_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_107_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_107_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_107_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_107_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_108_clock; // @[pe.scala 187:13]
  wire  PE_108_reset; // @[pe.scala 187:13]
  wire  PE_108_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_108_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_108_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_108_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_108_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_108_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_108_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_108_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_108_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_108_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_108_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_109_clock; // @[pe.scala 187:13]
  wire  PE_109_reset; // @[pe.scala 187:13]
  wire  PE_109_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_109_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_109_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_109_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_109_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_109_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_109_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_109_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_109_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_109_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_109_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_110_clock; // @[pe.scala 187:13]
  wire  PE_110_reset; // @[pe.scala 187:13]
  wire  PE_110_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_110_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_110_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_110_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_110_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_110_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_110_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_110_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_110_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_110_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_110_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_111_clock; // @[pe.scala 187:13]
  wire  PE_111_reset; // @[pe.scala 187:13]
  wire  PE_111_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_111_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_111_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_111_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_111_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_111_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_111_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_111_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_111_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_111_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_111_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_112_clock; // @[pe.scala 187:13]
  wire  PE_112_reset; // @[pe.scala 187:13]
  wire  PE_112_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_112_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_112_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_112_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_112_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_112_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_112_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_112_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_112_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_112_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_112_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_113_clock; // @[pe.scala 187:13]
  wire  PE_113_reset; // @[pe.scala 187:13]
  wire  PE_113_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_113_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_113_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_113_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_113_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_113_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_113_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_113_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_113_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_113_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_113_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_114_clock; // @[pe.scala 187:13]
  wire  PE_114_reset; // @[pe.scala 187:13]
  wire  PE_114_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_114_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_114_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_114_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_114_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_114_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_114_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_114_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_114_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_114_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_114_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_115_clock; // @[pe.scala 187:13]
  wire  PE_115_reset; // @[pe.scala 187:13]
  wire  PE_115_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_115_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_115_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_115_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_115_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_115_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_115_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_115_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_115_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_115_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_115_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_116_clock; // @[pe.scala 187:13]
  wire  PE_116_reset; // @[pe.scala 187:13]
  wire  PE_116_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_116_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_116_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_116_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_116_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_116_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_116_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_116_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_116_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_116_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_116_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_117_clock; // @[pe.scala 187:13]
  wire  PE_117_reset; // @[pe.scala 187:13]
  wire  PE_117_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_117_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_117_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_117_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_117_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_117_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_117_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_117_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_117_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_117_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_117_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_118_clock; // @[pe.scala 187:13]
  wire  PE_118_reset; // @[pe.scala 187:13]
  wire  PE_118_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_118_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_118_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_118_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_118_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_118_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_118_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_118_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_118_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_118_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_118_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_119_clock; // @[pe.scala 187:13]
  wire  PE_119_reset; // @[pe.scala 187:13]
  wire  PE_119_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_119_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_119_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_119_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_119_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_119_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_119_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_119_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_119_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_119_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_119_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_120_clock; // @[pe.scala 187:13]
  wire  PE_120_reset; // @[pe.scala 187:13]
  wire  PE_120_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_120_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_120_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_120_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_120_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_120_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_120_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_120_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_120_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_120_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_120_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_121_clock; // @[pe.scala 187:13]
  wire  PE_121_reset; // @[pe.scala 187:13]
  wire  PE_121_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_121_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_121_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_121_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_121_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_121_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_121_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_121_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_121_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_121_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_121_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_122_clock; // @[pe.scala 187:13]
  wire  PE_122_reset; // @[pe.scala 187:13]
  wire  PE_122_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_122_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_122_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_122_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_122_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_122_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_122_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_122_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_122_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_122_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_122_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_123_clock; // @[pe.scala 187:13]
  wire  PE_123_reset; // @[pe.scala 187:13]
  wire  PE_123_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_123_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_123_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_123_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_123_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_123_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_123_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_123_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_123_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_123_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_123_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_124_clock; // @[pe.scala 187:13]
  wire  PE_124_reset; // @[pe.scala 187:13]
  wire  PE_124_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_124_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_124_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_124_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_124_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_124_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_124_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_124_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_124_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_124_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_124_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_125_clock; // @[pe.scala 187:13]
  wire  PE_125_reset; // @[pe.scala 187:13]
  wire  PE_125_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_125_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_125_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_125_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_125_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_125_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_125_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_125_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_125_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_125_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_125_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_126_clock; // @[pe.scala 187:13]
  wire  PE_126_reset; // @[pe.scala 187:13]
  wire  PE_126_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_126_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_126_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_126_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_126_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_126_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_126_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_126_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_126_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_126_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_126_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_127_clock; // @[pe.scala 187:13]
  wire  PE_127_reset; // @[pe.scala 187:13]
  wire  PE_127_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_127_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_127_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_127_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_127_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_127_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_127_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_127_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_127_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_127_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_127_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_128_clock; // @[pe.scala 187:13]
  wire  PE_128_reset; // @[pe.scala 187:13]
  wire  PE_128_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_128_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_128_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_128_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_128_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_128_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_128_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_128_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_128_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_128_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_128_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_129_clock; // @[pe.scala 187:13]
  wire  PE_129_reset; // @[pe.scala 187:13]
  wire  PE_129_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_129_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_129_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_129_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_129_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_129_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_129_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_129_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_129_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_129_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_129_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_130_clock; // @[pe.scala 187:13]
  wire  PE_130_reset; // @[pe.scala 187:13]
  wire  PE_130_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_130_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_130_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_130_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_130_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_130_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_130_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_130_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_130_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_130_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_130_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_131_clock; // @[pe.scala 187:13]
  wire  PE_131_reset; // @[pe.scala 187:13]
  wire  PE_131_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_131_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_131_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_131_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_131_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_131_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_131_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_131_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_131_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_131_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_131_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_132_clock; // @[pe.scala 187:13]
  wire  PE_132_reset; // @[pe.scala 187:13]
  wire  PE_132_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_132_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_132_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_132_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_132_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_132_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_132_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_132_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_132_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_132_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_132_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_133_clock; // @[pe.scala 187:13]
  wire  PE_133_reset; // @[pe.scala 187:13]
  wire  PE_133_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_133_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_133_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_133_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_133_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_133_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_133_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_133_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_133_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_133_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_133_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_134_clock; // @[pe.scala 187:13]
  wire  PE_134_reset; // @[pe.scala 187:13]
  wire  PE_134_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_134_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_134_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_134_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_134_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_134_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_134_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_134_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_134_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_134_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_134_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_135_clock; // @[pe.scala 187:13]
  wire  PE_135_reset; // @[pe.scala 187:13]
  wire  PE_135_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_135_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_135_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_135_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_135_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_135_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_135_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_135_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_135_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_135_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_135_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_136_clock; // @[pe.scala 187:13]
  wire  PE_136_reset; // @[pe.scala 187:13]
  wire  PE_136_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_136_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_136_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_136_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_136_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_136_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_136_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_136_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_136_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_136_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_136_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_137_clock; // @[pe.scala 187:13]
  wire  PE_137_reset; // @[pe.scala 187:13]
  wire  PE_137_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_137_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_137_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_137_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_137_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_137_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_137_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_137_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_137_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_137_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_137_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_138_clock; // @[pe.scala 187:13]
  wire  PE_138_reset; // @[pe.scala 187:13]
  wire  PE_138_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_138_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_138_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_138_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_138_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_138_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_138_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_138_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_138_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_138_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_138_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_139_clock; // @[pe.scala 187:13]
  wire  PE_139_reset; // @[pe.scala 187:13]
  wire  PE_139_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_139_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_139_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_139_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_139_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_139_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_139_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_139_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_139_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_139_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_139_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_140_clock; // @[pe.scala 187:13]
  wire  PE_140_reset; // @[pe.scala 187:13]
  wire  PE_140_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_140_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_140_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_140_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_140_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_140_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_140_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_140_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_140_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_140_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_140_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_141_clock; // @[pe.scala 187:13]
  wire  PE_141_reset; // @[pe.scala 187:13]
  wire  PE_141_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_141_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_141_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_141_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_141_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_141_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_141_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_141_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_141_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_141_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_141_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_142_clock; // @[pe.scala 187:13]
  wire  PE_142_reset; // @[pe.scala 187:13]
  wire  PE_142_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_142_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_142_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_142_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_142_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_142_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_142_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_142_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_142_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_142_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_142_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_143_clock; // @[pe.scala 187:13]
  wire  PE_143_reset; // @[pe.scala 187:13]
  wire  PE_143_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_143_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_143_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_143_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_143_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_143_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_143_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_143_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_143_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_143_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_143_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_144_clock; // @[pe.scala 187:13]
  wire  PE_144_reset; // @[pe.scala 187:13]
  wire  PE_144_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_144_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_144_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_144_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_144_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_144_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_144_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_144_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_144_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_144_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_144_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_145_clock; // @[pe.scala 187:13]
  wire  PE_145_reset; // @[pe.scala 187:13]
  wire  PE_145_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_145_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_145_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_145_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_145_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_145_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_145_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_145_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_145_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_145_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_145_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_146_clock; // @[pe.scala 187:13]
  wire  PE_146_reset; // @[pe.scala 187:13]
  wire  PE_146_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_146_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_146_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_146_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_146_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_146_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_146_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_146_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_146_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_146_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_146_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_147_clock; // @[pe.scala 187:13]
  wire  PE_147_reset; // @[pe.scala 187:13]
  wire  PE_147_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_147_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_147_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_147_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_147_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_147_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_147_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_147_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_147_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_147_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_147_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_148_clock; // @[pe.scala 187:13]
  wire  PE_148_reset; // @[pe.scala 187:13]
  wire  PE_148_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_148_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_148_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_148_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_148_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_148_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_148_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_148_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_148_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_148_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_148_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_149_clock; // @[pe.scala 187:13]
  wire  PE_149_reset; // @[pe.scala 187:13]
  wire  PE_149_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_149_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_149_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_149_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_149_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_149_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_149_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_149_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_149_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_149_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_149_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_150_clock; // @[pe.scala 187:13]
  wire  PE_150_reset; // @[pe.scala 187:13]
  wire  PE_150_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_150_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_150_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_150_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_150_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_150_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_150_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_150_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_150_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_150_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_150_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_151_clock; // @[pe.scala 187:13]
  wire  PE_151_reset; // @[pe.scala 187:13]
  wire  PE_151_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_151_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_151_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_151_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_151_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_151_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_151_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_151_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_151_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_151_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_151_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_152_clock; // @[pe.scala 187:13]
  wire  PE_152_reset; // @[pe.scala 187:13]
  wire  PE_152_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_152_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_152_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_152_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_152_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_152_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_152_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_152_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_152_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_152_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_152_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_153_clock; // @[pe.scala 187:13]
  wire  PE_153_reset; // @[pe.scala 187:13]
  wire  PE_153_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_153_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_153_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_153_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_153_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_153_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_153_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_153_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_153_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_153_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_153_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_154_clock; // @[pe.scala 187:13]
  wire  PE_154_reset; // @[pe.scala 187:13]
  wire  PE_154_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_154_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_154_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_154_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_154_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_154_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_154_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_154_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_154_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_154_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_154_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_155_clock; // @[pe.scala 187:13]
  wire  PE_155_reset; // @[pe.scala 187:13]
  wire  PE_155_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_155_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_155_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_155_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_155_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_155_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_155_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_155_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_155_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_155_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_155_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_156_clock; // @[pe.scala 187:13]
  wire  PE_156_reset; // @[pe.scala 187:13]
  wire  PE_156_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_156_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_156_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_156_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_156_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_156_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_156_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_156_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_156_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_156_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_156_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_157_clock; // @[pe.scala 187:13]
  wire  PE_157_reset; // @[pe.scala 187:13]
  wire  PE_157_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_157_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_157_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_157_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_157_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_157_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_157_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_157_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_157_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_157_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_157_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_158_clock; // @[pe.scala 187:13]
  wire  PE_158_reset; // @[pe.scala 187:13]
  wire  PE_158_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_158_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_158_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_158_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_158_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_158_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_158_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_158_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_158_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_158_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_158_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_159_clock; // @[pe.scala 187:13]
  wire  PE_159_reset; // @[pe.scala 187:13]
  wire  PE_159_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_159_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_159_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_159_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_159_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_159_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_159_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_159_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_159_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_159_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_159_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_160_clock; // @[pe.scala 187:13]
  wire  PE_160_reset; // @[pe.scala 187:13]
  wire  PE_160_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_160_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_160_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_160_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_160_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_160_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_160_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_160_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_160_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_160_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_160_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_161_clock; // @[pe.scala 187:13]
  wire  PE_161_reset; // @[pe.scala 187:13]
  wire  PE_161_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_161_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_161_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_161_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_161_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_161_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_161_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_161_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_161_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_161_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_161_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_162_clock; // @[pe.scala 187:13]
  wire  PE_162_reset; // @[pe.scala 187:13]
  wire  PE_162_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_162_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_162_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_162_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_162_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_162_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_162_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_162_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_162_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_162_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_162_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_163_clock; // @[pe.scala 187:13]
  wire  PE_163_reset; // @[pe.scala 187:13]
  wire  PE_163_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_163_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_163_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_163_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_163_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_163_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_163_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_163_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_163_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_163_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_163_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_164_clock; // @[pe.scala 187:13]
  wire  PE_164_reset; // @[pe.scala 187:13]
  wire  PE_164_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_164_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_164_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_164_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_164_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_164_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_164_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_164_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_164_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_164_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_164_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_165_clock; // @[pe.scala 187:13]
  wire  PE_165_reset; // @[pe.scala 187:13]
  wire  PE_165_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_165_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_165_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_165_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_165_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_165_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_165_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_165_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_165_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_165_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_165_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_166_clock; // @[pe.scala 187:13]
  wire  PE_166_reset; // @[pe.scala 187:13]
  wire  PE_166_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_166_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_166_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_166_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_166_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_166_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_166_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_166_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_166_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_166_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_166_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_167_clock; // @[pe.scala 187:13]
  wire  PE_167_reset; // @[pe.scala 187:13]
  wire  PE_167_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_167_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_167_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_167_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_167_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_167_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_167_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_167_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_167_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_167_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_167_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_168_clock; // @[pe.scala 187:13]
  wire  PE_168_reset; // @[pe.scala 187:13]
  wire  PE_168_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_168_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_168_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_168_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_168_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_168_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_168_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_168_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_168_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_168_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_168_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_169_clock; // @[pe.scala 187:13]
  wire  PE_169_reset; // @[pe.scala 187:13]
  wire  PE_169_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_169_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_169_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_169_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_169_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_169_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_169_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_169_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_169_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_169_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_169_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_170_clock; // @[pe.scala 187:13]
  wire  PE_170_reset; // @[pe.scala 187:13]
  wire  PE_170_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_170_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_170_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_170_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_170_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_170_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_170_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_170_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_170_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_170_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_170_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_171_clock; // @[pe.scala 187:13]
  wire  PE_171_reset; // @[pe.scala 187:13]
  wire  PE_171_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_171_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_171_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_171_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_171_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_171_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_171_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_171_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_171_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_171_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_171_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_172_clock; // @[pe.scala 187:13]
  wire  PE_172_reset; // @[pe.scala 187:13]
  wire  PE_172_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_172_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_172_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_172_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_172_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_172_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_172_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_172_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_172_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_172_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_172_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_173_clock; // @[pe.scala 187:13]
  wire  PE_173_reset; // @[pe.scala 187:13]
  wire  PE_173_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_173_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_173_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_173_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_173_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_173_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_173_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_173_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_173_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_173_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_173_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_174_clock; // @[pe.scala 187:13]
  wire  PE_174_reset; // @[pe.scala 187:13]
  wire  PE_174_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_174_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_174_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_174_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_174_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_174_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_174_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_174_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_174_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_174_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_174_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_175_clock; // @[pe.scala 187:13]
  wire  PE_175_reset; // @[pe.scala 187:13]
  wire  PE_175_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_175_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_175_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_175_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_175_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_175_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_175_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_175_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_175_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_175_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_175_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_176_clock; // @[pe.scala 187:13]
  wire  PE_176_reset; // @[pe.scala 187:13]
  wire  PE_176_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_176_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_176_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_176_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_176_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_176_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_176_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_176_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_176_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_176_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_176_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_177_clock; // @[pe.scala 187:13]
  wire  PE_177_reset; // @[pe.scala 187:13]
  wire  PE_177_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_177_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_177_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_177_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_177_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_177_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_177_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_177_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_177_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_177_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_177_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_178_clock; // @[pe.scala 187:13]
  wire  PE_178_reset; // @[pe.scala 187:13]
  wire  PE_178_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_178_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_178_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_178_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_178_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_178_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_178_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_178_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_178_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_178_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_178_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_179_clock; // @[pe.scala 187:13]
  wire  PE_179_reset; // @[pe.scala 187:13]
  wire  PE_179_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_179_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_179_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_179_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_179_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_179_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_179_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_179_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_179_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_179_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_179_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_180_clock; // @[pe.scala 187:13]
  wire  PE_180_reset; // @[pe.scala 187:13]
  wire  PE_180_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_180_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_180_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_180_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_180_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_180_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_180_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_180_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_180_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_180_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_180_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_181_clock; // @[pe.scala 187:13]
  wire  PE_181_reset; // @[pe.scala 187:13]
  wire  PE_181_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_181_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_181_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_181_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_181_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_181_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_181_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_181_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_181_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_181_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_181_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_182_clock; // @[pe.scala 187:13]
  wire  PE_182_reset; // @[pe.scala 187:13]
  wire  PE_182_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_182_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_182_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_182_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_182_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_182_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_182_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_182_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_182_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_182_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_182_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_183_clock; // @[pe.scala 187:13]
  wire  PE_183_reset; // @[pe.scala 187:13]
  wire  PE_183_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_183_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_183_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_183_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_183_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_183_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_183_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_183_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_183_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_183_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_183_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_184_clock; // @[pe.scala 187:13]
  wire  PE_184_reset; // @[pe.scala 187:13]
  wire  PE_184_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_184_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_184_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_184_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_184_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_184_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_184_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_184_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_184_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_184_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_184_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_185_clock; // @[pe.scala 187:13]
  wire  PE_185_reset; // @[pe.scala 187:13]
  wire  PE_185_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_185_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_185_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_185_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_185_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_185_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_185_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_185_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_185_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_185_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_185_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_186_clock; // @[pe.scala 187:13]
  wire  PE_186_reset; // @[pe.scala 187:13]
  wire  PE_186_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_186_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_186_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_186_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_186_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_186_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_186_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_186_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_186_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_186_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_186_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_187_clock; // @[pe.scala 187:13]
  wire  PE_187_reset; // @[pe.scala 187:13]
  wire  PE_187_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_187_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_187_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_187_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_187_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_187_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_187_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_187_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_187_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_187_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_187_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_188_clock; // @[pe.scala 187:13]
  wire  PE_188_reset; // @[pe.scala 187:13]
  wire  PE_188_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_188_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_188_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_188_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_188_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_188_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_188_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_188_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_188_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_188_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_188_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_189_clock; // @[pe.scala 187:13]
  wire  PE_189_reset; // @[pe.scala 187:13]
  wire  PE_189_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_189_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_189_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_189_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_189_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_189_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_189_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_189_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_189_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_189_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_189_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_190_clock; // @[pe.scala 187:13]
  wire  PE_190_reset; // @[pe.scala 187:13]
  wire  PE_190_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_190_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_190_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_190_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_190_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_190_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_190_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_190_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_190_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_190_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_190_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_191_clock; // @[pe.scala 187:13]
  wire  PE_191_reset; // @[pe.scala 187:13]
  wire  PE_191_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_191_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_191_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_191_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_191_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_191_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_191_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_191_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_191_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_191_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_191_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_192_clock; // @[pe.scala 187:13]
  wire  PE_192_reset; // @[pe.scala 187:13]
  wire  PE_192_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_192_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_192_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_192_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_192_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_192_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_192_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_192_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_192_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_192_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_192_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_193_clock; // @[pe.scala 187:13]
  wire  PE_193_reset; // @[pe.scala 187:13]
  wire  PE_193_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_193_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_193_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_193_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_193_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_193_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_193_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_193_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_193_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_193_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_193_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_194_clock; // @[pe.scala 187:13]
  wire  PE_194_reset; // @[pe.scala 187:13]
  wire  PE_194_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_194_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_194_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_194_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_194_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_194_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_194_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_194_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_194_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_194_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_194_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_195_clock; // @[pe.scala 187:13]
  wire  PE_195_reset; // @[pe.scala 187:13]
  wire  PE_195_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_195_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_195_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_195_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_195_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_195_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_195_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_195_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_195_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_195_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_195_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_196_clock; // @[pe.scala 187:13]
  wire  PE_196_reset; // @[pe.scala 187:13]
  wire  PE_196_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_196_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_196_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_196_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_196_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_196_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_196_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_196_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_196_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_196_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_196_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_197_clock; // @[pe.scala 187:13]
  wire  PE_197_reset; // @[pe.scala 187:13]
  wire  PE_197_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_197_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_197_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_197_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_197_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_197_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_197_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_197_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_197_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_197_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_197_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_198_clock; // @[pe.scala 187:13]
  wire  PE_198_reset; // @[pe.scala 187:13]
  wire  PE_198_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_198_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_198_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_198_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_198_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_198_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_198_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_198_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_198_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_198_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_198_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_199_clock; // @[pe.scala 187:13]
  wire  PE_199_reset; // @[pe.scala 187:13]
  wire  PE_199_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_199_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_199_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_199_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_199_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_199_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_199_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_199_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_199_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_199_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_199_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_200_clock; // @[pe.scala 187:13]
  wire  PE_200_reset; // @[pe.scala 187:13]
  wire  PE_200_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_200_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_200_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_200_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_200_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_200_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_200_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_200_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_200_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_200_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_200_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_201_clock; // @[pe.scala 187:13]
  wire  PE_201_reset; // @[pe.scala 187:13]
  wire  PE_201_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_201_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_201_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_201_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_201_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_201_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_201_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_201_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_201_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_201_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_201_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_202_clock; // @[pe.scala 187:13]
  wire  PE_202_reset; // @[pe.scala 187:13]
  wire  PE_202_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_202_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_202_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_202_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_202_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_202_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_202_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_202_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_202_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_202_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_202_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_203_clock; // @[pe.scala 187:13]
  wire  PE_203_reset; // @[pe.scala 187:13]
  wire  PE_203_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_203_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_203_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_203_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_203_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_203_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_203_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_203_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_203_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_203_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_203_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_204_clock; // @[pe.scala 187:13]
  wire  PE_204_reset; // @[pe.scala 187:13]
  wire  PE_204_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_204_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_204_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_204_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_204_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_204_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_204_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_204_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_204_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_204_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_204_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_205_clock; // @[pe.scala 187:13]
  wire  PE_205_reset; // @[pe.scala 187:13]
  wire  PE_205_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_205_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_205_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_205_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_205_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_205_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_205_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_205_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_205_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_205_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_205_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_206_clock; // @[pe.scala 187:13]
  wire  PE_206_reset; // @[pe.scala 187:13]
  wire  PE_206_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_206_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_206_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_206_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_206_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_206_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_206_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_206_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_206_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_206_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_206_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_207_clock; // @[pe.scala 187:13]
  wire  PE_207_reset; // @[pe.scala 187:13]
  wire  PE_207_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_207_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_207_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_207_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_207_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_207_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_207_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_207_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_207_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_207_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_207_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_208_clock; // @[pe.scala 187:13]
  wire  PE_208_reset; // @[pe.scala 187:13]
  wire  PE_208_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_208_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_208_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_208_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_208_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_208_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_208_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_208_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_208_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_208_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_208_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_209_clock; // @[pe.scala 187:13]
  wire  PE_209_reset; // @[pe.scala 187:13]
  wire  PE_209_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_209_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_209_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_209_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_209_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_209_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_209_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_209_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_209_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_209_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_209_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_210_clock; // @[pe.scala 187:13]
  wire  PE_210_reset; // @[pe.scala 187:13]
  wire  PE_210_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_210_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_210_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_210_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_210_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_210_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_210_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_210_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_210_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_210_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_210_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_211_clock; // @[pe.scala 187:13]
  wire  PE_211_reset; // @[pe.scala 187:13]
  wire  PE_211_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_211_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_211_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_211_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_211_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_211_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_211_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_211_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_211_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_211_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_211_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_212_clock; // @[pe.scala 187:13]
  wire  PE_212_reset; // @[pe.scala 187:13]
  wire  PE_212_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_212_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_212_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_212_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_212_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_212_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_212_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_212_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_212_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_212_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_212_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_213_clock; // @[pe.scala 187:13]
  wire  PE_213_reset; // @[pe.scala 187:13]
  wire  PE_213_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_213_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_213_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_213_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_213_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_213_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_213_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_213_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_213_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_213_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_213_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_214_clock; // @[pe.scala 187:13]
  wire  PE_214_reset; // @[pe.scala 187:13]
  wire  PE_214_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_214_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_214_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_214_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_214_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_214_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_214_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_214_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_214_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_214_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_214_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_215_clock; // @[pe.scala 187:13]
  wire  PE_215_reset; // @[pe.scala 187:13]
  wire  PE_215_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_215_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_215_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_215_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_215_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_215_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_215_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_215_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_215_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_215_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_215_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_216_clock; // @[pe.scala 187:13]
  wire  PE_216_reset; // @[pe.scala 187:13]
  wire  PE_216_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_216_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_216_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_216_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_216_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_216_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_216_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_216_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_216_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_216_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_216_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_217_clock; // @[pe.scala 187:13]
  wire  PE_217_reset; // @[pe.scala 187:13]
  wire  PE_217_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_217_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_217_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_217_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_217_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_217_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_217_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_217_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_217_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_217_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_217_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_218_clock; // @[pe.scala 187:13]
  wire  PE_218_reset; // @[pe.scala 187:13]
  wire  PE_218_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_218_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_218_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_218_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_218_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_218_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_218_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_218_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_218_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_218_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_218_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_219_clock; // @[pe.scala 187:13]
  wire  PE_219_reset; // @[pe.scala 187:13]
  wire  PE_219_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_219_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_219_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_219_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_219_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_219_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_219_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_219_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_219_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_219_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_219_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_220_clock; // @[pe.scala 187:13]
  wire  PE_220_reset; // @[pe.scala 187:13]
  wire  PE_220_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_220_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_220_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_220_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_220_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_220_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_220_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_220_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_220_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_220_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_220_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_221_clock; // @[pe.scala 187:13]
  wire  PE_221_reset; // @[pe.scala 187:13]
  wire  PE_221_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_221_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_221_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_221_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_221_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_221_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_221_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_221_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_221_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_221_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_221_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_222_clock; // @[pe.scala 187:13]
  wire  PE_222_reset; // @[pe.scala 187:13]
  wire  PE_222_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_222_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_222_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_222_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_222_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_222_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_222_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_222_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_222_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_222_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_222_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_223_clock; // @[pe.scala 187:13]
  wire  PE_223_reset; // @[pe.scala 187:13]
  wire  PE_223_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_223_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_223_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_223_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_223_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_223_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_223_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_223_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_223_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_223_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_223_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_224_clock; // @[pe.scala 187:13]
  wire  PE_224_reset; // @[pe.scala 187:13]
  wire  PE_224_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_224_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_224_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_224_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_224_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_224_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_224_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_224_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_224_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_224_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_224_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_225_clock; // @[pe.scala 187:13]
  wire  PE_225_reset; // @[pe.scala 187:13]
  wire  PE_225_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_225_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_225_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_225_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_225_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_225_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_225_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_225_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_225_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_225_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_225_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_226_clock; // @[pe.scala 187:13]
  wire  PE_226_reset; // @[pe.scala 187:13]
  wire  PE_226_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_226_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_226_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_226_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_226_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_226_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_226_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_226_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_226_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_226_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_226_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_227_clock; // @[pe.scala 187:13]
  wire  PE_227_reset; // @[pe.scala 187:13]
  wire  PE_227_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_227_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_227_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_227_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_227_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_227_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_227_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_227_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_227_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_227_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_227_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_228_clock; // @[pe.scala 187:13]
  wire  PE_228_reset; // @[pe.scala 187:13]
  wire  PE_228_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_228_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_228_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_228_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_228_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_228_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_228_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_228_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_228_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_228_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_228_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_229_clock; // @[pe.scala 187:13]
  wire  PE_229_reset; // @[pe.scala 187:13]
  wire  PE_229_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_229_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_229_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_229_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_229_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_229_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_229_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_229_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_229_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_229_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_229_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_230_clock; // @[pe.scala 187:13]
  wire  PE_230_reset; // @[pe.scala 187:13]
  wire  PE_230_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_230_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_230_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_230_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_230_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_230_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_230_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_230_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_230_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_230_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_230_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_231_clock; // @[pe.scala 187:13]
  wire  PE_231_reset; // @[pe.scala 187:13]
  wire  PE_231_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_231_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_231_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_231_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_231_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_231_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_231_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_231_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_231_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_231_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_231_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_232_clock; // @[pe.scala 187:13]
  wire  PE_232_reset; // @[pe.scala 187:13]
  wire  PE_232_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_232_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_232_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_232_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_232_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_232_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_232_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_232_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_232_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_232_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_232_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_233_clock; // @[pe.scala 187:13]
  wire  PE_233_reset; // @[pe.scala 187:13]
  wire  PE_233_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_233_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_233_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_233_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_233_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_233_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_233_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_233_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_233_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_233_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_233_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_234_clock; // @[pe.scala 187:13]
  wire  PE_234_reset; // @[pe.scala 187:13]
  wire  PE_234_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_234_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_234_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_234_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_234_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_234_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_234_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_234_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_234_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_234_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_234_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_235_clock; // @[pe.scala 187:13]
  wire  PE_235_reset; // @[pe.scala 187:13]
  wire  PE_235_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_235_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_235_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_235_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_235_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_235_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_235_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_235_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_235_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_235_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_235_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_236_clock; // @[pe.scala 187:13]
  wire  PE_236_reset; // @[pe.scala 187:13]
  wire  PE_236_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_236_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_236_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_236_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_236_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_236_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_236_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_236_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_236_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_236_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_236_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_237_clock; // @[pe.scala 187:13]
  wire  PE_237_reset; // @[pe.scala 187:13]
  wire  PE_237_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_237_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_237_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_237_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_237_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_237_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_237_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_237_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_237_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_237_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_237_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_238_clock; // @[pe.scala 187:13]
  wire  PE_238_reset; // @[pe.scala 187:13]
  wire  PE_238_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_238_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_238_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_238_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_238_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_238_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_238_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_238_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_238_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_238_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_238_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_239_clock; // @[pe.scala 187:13]
  wire  PE_239_reset; // @[pe.scala 187:13]
  wire  PE_239_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_239_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_239_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_239_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_239_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_239_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_239_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_239_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_239_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_239_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_239_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_240_clock; // @[pe.scala 187:13]
  wire  PE_240_reset; // @[pe.scala 187:13]
  wire  PE_240_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_240_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_240_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_240_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_240_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_240_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_240_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_240_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_240_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_240_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_240_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_241_clock; // @[pe.scala 187:13]
  wire  PE_241_reset; // @[pe.scala 187:13]
  wire  PE_241_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_241_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_241_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_241_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_241_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_241_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_241_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_241_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_241_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_241_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_241_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_242_clock; // @[pe.scala 187:13]
  wire  PE_242_reset; // @[pe.scala 187:13]
  wire  PE_242_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_242_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_242_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_242_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_242_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_242_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_242_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_242_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_242_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_242_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_242_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_243_clock; // @[pe.scala 187:13]
  wire  PE_243_reset; // @[pe.scala 187:13]
  wire  PE_243_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_243_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_243_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_243_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_243_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_243_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_243_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_243_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_243_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_243_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_243_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_244_clock; // @[pe.scala 187:13]
  wire  PE_244_reset; // @[pe.scala 187:13]
  wire  PE_244_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_244_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_244_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_244_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_244_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_244_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_244_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_244_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_244_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_244_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_244_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_245_clock; // @[pe.scala 187:13]
  wire  PE_245_reset; // @[pe.scala 187:13]
  wire  PE_245_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_245_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_245_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_245_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_245_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_245_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_245_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_245_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_245_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_245_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_245_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_246_clock; // @[pe.scala 187:13]
  wire  PE_246_reset; // @[pe.scala 187:13]
  wire  PE_246_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_246_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_246_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_246_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_246_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_246_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_246_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_246_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_246_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_246_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_246_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_247_clock; // @[pe.scala 187:13]
  wire  PE_247_reset; // @[pe.scala 187:13]
  wire  PE_247_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_247_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_247_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_247_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_247_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_247_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_247_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_247_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_247_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_247_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_247_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_248_clock; // @[pe.scala 187:13]
  wire  PE_248_reset; // @[pe.scala 187:13]
  wire  PE_248_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_248_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_248_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_248_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_248_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_248_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_248_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_248_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_248_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_248_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_248_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_249_clock; // @[pe.scala 187:13]
  wire  PE_249_reset; // @[pe.scala 187:13]
  wire  PE_249_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_249_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_249_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_249_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_249_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_249_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_249_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_249_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_249_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_249_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_249_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_250_clock; // @[pe.scala 187:13]
  wire  PE_250_reset; // @[pe.scala 187:13]
  wire  PE_250_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_250_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_250_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_250_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_250_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_250_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_250_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_250_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_250_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_250_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_250_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_251_clock; // @[pe.scala 187:13]
  wire  PE_251_reset; // @[pe.scala 187:13]
  wire  PE_251_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_251_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_251_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_251_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_251_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_251_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_251_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_251_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_251_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_251_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_251_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_252_clock; // @[pe.scala 187:13]
  wire  PE_252_reset; // @[pe.scala 187:13]
  wire  PE_252_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_252_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_252_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_252_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_252_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_252_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_252_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_252_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_252_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_252_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_252_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_253_clock; // @[pe.scala 187:13]
  wire  PE_253_reset; // @[pe.scala 187:13]
  wire  PE_253_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_253_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_253_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_253_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_253_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_253_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_253_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_253_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_253_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_253_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_253_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_254_clock; // @[pe.scala 187:13]
  wire  PE_254_reset; // @[pe.scala 187:13]
  wire  PE_254_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_254_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_254_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_254_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_254_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_254_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_254_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_254_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_254_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_254_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_254_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_255_clock; // @[pe.scala 187:13]
  wire  PE_255_reset; // @[pe.scala 187:13]
  wire  PE_255_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_255_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_255_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_255_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_255_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_255_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_255_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_255_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_255_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_255_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_255_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_256_clock; // @[pe.scala 187:13]
  wire  PE_256_reset; // @[pe.scala 187:13]
  wire  PE_256_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_256_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_256_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_256_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_256_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_256_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_256_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_256_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_256_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_256_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_256_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_257_clock; // @[pe.scala 187:13]
  wire  PE_257_reset; // @[pe.scala 187:13]
  wire  PE_257_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_257_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_257_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_257_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_257_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_257_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_257_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_257_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_257_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_257_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_257_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_258_clock; // @[pe.scala 187:13]
  wire  PE_258_reset; // @[pe.scala 187:13]
  wire  PE_258_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_258_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_258_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_258_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_258_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_258_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_258_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_258_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_258_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_258_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_258_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_259_clock; // @[pe.scala 187:13]
  wire  PE_259_reset; // @[pe.scala 187:13]
  wire  PE_259_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_259_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_259_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_259_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_259_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_259_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_259_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_259_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_259_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_259_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_259_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_260_clock; // @[pe.scala 187:13]
  wire  PE_260_reset; // @[pe.scala 187:13]
  wire  PE_260_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_260_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_260_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_260_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_260_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_260_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_260_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_260_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_260_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_260_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_260_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_261_clock; // @[pe.scala 187:13]
  wire  PE_261_reset; // @[pe.scala 187:13]
  wire  PE_261_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_261_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_261_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_261_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_261_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_261_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_261_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_261_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_261_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_261_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_261_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_262_clock; // @[pe.scala 187:13]
  wire  PE_262_reset; // @[pe.scala 187:13]
  wire  PE_262_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_262_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_262_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_262_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_262_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_262_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_262_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_262_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_262_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_262_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_262_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_263_clock; // @[pe.scala 187:13]
  wire  PE_263_reset; // @[pe.scala 187:13]
  wire  PE_263_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_263_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_263_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_263_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_263_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_263_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_263_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_263_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_263_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_263_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_263_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_264_clock; // @[pe.scala 187:13]
  wire  PE_264_reset; // @[pe.scala 187:13]
  wire  PE_264_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_264_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_264_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_264_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_264_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_264_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_264_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_264_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_264_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_264_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_264_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_265_clock; // @[pe.scala 187:13]
  wire  PE_265_reset; // @[pe.scala 187:13]
  wire  PE_265_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_265_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_265_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_265_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_265_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_265_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_265_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_265_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_265_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_265_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_265_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_266_clock; // @[pe.scala 187:13]
  wire  PE_266_reset; // @[pe.scala 187:13]
  wire  PE_266_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_266_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_266_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_266_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_266_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_266_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_266_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_266_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_266_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_266_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_266_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_267_clock; // @[pe.scala 187:13]
  wire  PE_267_reset; // @[pe.scala 187:13]
  wire  PE_267_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_267_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_267_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_267_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_267_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_267_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_267_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_267_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_267_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_267_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_267_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_268_clock; // @[pe.scala 187:13]
  wire  PE_268_reset; // @[pe.scala 187:13]
  wire  PE_268_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_268_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_268_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_268_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_268_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_268_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_268_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_268_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_268_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_268_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_268_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_269_clock; // @[pe.scala 187:13]
  wire  PE_269_reset; // @[pe.scala 187:13]
  wire  PE_269_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_269_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_269_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_269_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_269_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_269_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_269_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_269_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_269_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_269_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_269_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_270_clock; // @[pe.scala 187:13]
  wire  PE_270_reset; // @[pe.scala 187:13]
  wire  PE_270_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_270_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_270_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_270_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_270_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_270_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_270_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_270_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_270_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_270_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_270_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_271_clock; // @[pe.scala 187:13]
  wire  PE_271_reset; // @[pe.scala 187:13]
  wire  PE_271_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_271_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_271_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_271_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_271_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_271_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_271_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_271_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_271_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_271_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_271_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_272_clock; // @[pe.scala 187:13]
  wire  PE_272_reset; // @[pe.scala 187:13]
  wire  PE_272_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_272_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_272_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_272_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_272_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_272_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_272_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_272_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_272_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_272_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_272_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_273_clock; // @[pe.scala 187:13]
  wire  PE_273_reset; // @[pe.scala 187:13]
  wire  PE_273_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_273_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_273_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_273_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_273_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_273_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_273_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_273_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_273_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_273_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_273_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_274_clock; // @[pe.scala 187:13]
  wire  PE_274_reset; // @[pe.scala 187:13]
  wire  PE_274_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_274_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_274_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_274_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_274_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_274_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_274_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_274_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_274_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_274_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_274_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_275_clock; // @[pe.scala 187:13]
  wire  PE_275_reset; // @[pe.scala 187:13]
  wire  PE_275_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_275_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_275_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_275_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_275_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_275_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_275_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_275_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_275_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_275_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_275_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_276_clock; // @[pe.scala 187:13]
  wire  PE_276_reset; // @[pe.scala 187:13]
  wire  PE_276_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_276_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_276_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_276_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_276_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_276_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_276_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_276_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_276_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_276_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_276_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_277_clock; // @[pe.scala 187:13]
  wire  PE_277_reset; // @[pe.scala 187:13]
  wire  PE_277_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_277_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_277_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_277_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_277_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_277_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_277_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_277_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_277_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_277_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_277_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_278_clock; // @[pe.scala 187:13]
  wire  PE_278_reset; // @[pe.scala 187:13]
  wire  PE_278_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_278_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_278_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_278_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_278_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_278_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_278_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_278_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_278_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_278_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_278_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_279_clock; // @[pe.scala 187:13]
  wire  PE_279_reset; // @[pe.scala 187:13]
  wire  PE_279_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_279_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_279_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_279_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_279_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_279_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_279_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_279_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_279_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_279_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_279_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_280_clock; // @[pe.scala 187:13]
  wire  PE_280_reset; // @[pe.scala 187:13]
  wire  PE_280_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_280_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_280_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_280_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_280_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_280_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_280_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_280_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_280_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_280_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_280_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_281_clock; // @[pe.scala 187:13]
  wire  PE_281_reset; // @[pe.scala 187:13]
  wire  PE_281_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_281_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_281_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_281_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_281_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_281_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_281_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_281_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_281_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_281_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_281_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_282_clock; // @[pe.scala 187:13]
  wire  PE_282_reset; // @[pe.scala 187:13]
  wire  PE_282_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_282_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_282_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_282_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_282_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_282_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_282_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_282_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_282_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_282_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_282_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_283_clock; // @[pe.scala 187:13]
  wire  PE_283_reset; // @[pe.scala 187:13]
  wire  PE_283_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_283_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_283_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_283_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_283_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_283_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_283_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_283_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_283_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_283_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_283_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_284_clock; // @[pe.scala 187:13]
  wire  PE_284_reset; // @[pe.scala 187:13]
  wire  PE_284_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_284_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_284_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_284_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_284_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_284_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_284_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_284_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_284_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_284_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_284_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_285_clock; // @[pe.scala 187:13]
  wire  PE_285_reset; // @[pe.scala 187:13]
  wire  PE_285_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_285_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_285_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_285_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_285_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_285_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_285_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_285_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_285_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_285_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_285_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_286_clock; // @[pe.scala 187:13]
  wire  PE_286_reset; // @[pe.scala 187:13]
  wire  PE_286_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_286_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_286_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_286_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_286_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_286_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_286_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_286_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_286_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_286_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_286_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_287_clock; // @[pe.scala 187:13]
  wire  PE_287_reset; // @[pe.scala 187:13]
  wire  PE_287_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_287_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_287_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_287_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_287_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_287_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_287_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_287_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_287_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_287_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_287_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_288_clock; // @[pe.scala 187:13]
  wire  PE_288_reset; // @[pe.scala 187:13]
  wire  PE_288_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_288_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_288_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_288_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_288_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_288_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_288_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_288_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_288_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_288_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_288_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_289_clock; // @[pe.scala 187:13]
  wire  PE_289_reset; // @[pe.scala 187:13]
  wire  PE_289_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_289_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_289_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_289_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_289_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_289_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_289_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_289_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_289_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_289_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_289_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_290_clock; // @[pe.scala 187:13]
  wire  PE_290_reset; // @[pe.scala 187:13]
  wire  PE_290_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_290_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_290_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_290_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_290_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_290_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_290_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_290_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_290_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_290_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_290_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_291_clock; // @[pe.scala 187:13]
  wire  PE_291_reset; // @[pe.scala 187:13]
  wire  PE_291_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_291_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_291_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_291_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_291_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_291_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_291_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_291_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_291_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_291_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_291_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_292_clock; // @[pe.scala 187:13]
  wire  PE_292_reset; // @[pe.scala 187:13]
  wire  PE_292_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_292_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_292_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_292_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_292_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_292_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_292_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_292_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_292_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_292_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_292_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_293_clock; // @[pe.scala 187:13]
  wire  PE_293_reset; // @[pe.scala 187:13]
  wire  PE_293_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_293_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_293_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_293_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_293_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_293_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_293_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_293_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_293_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_293_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_293_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_294_clock; // @[pe.scala 187:13]
  wire  PE_294_reset; // @[pe.scala 187:13]
  wire  PE_294_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_294_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_294_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_294_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_294_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_294_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_294_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_294_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_294_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_294_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_294_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_295_clock; // @[pe.scala 187:13]
  wire  PE_295_reset; // @[pe.scala 187:13]
  wire  PE_295_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_295_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_295_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_295_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_295_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_295_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_295_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_295_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_295_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_295_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_295_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_296_clock; // @[pe.scala 187:13]
  wire  PE_296_reset; // @[pe.scala 187:13]
  wire  PE_296_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_296_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_296_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_296_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_296_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_296_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_296_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_296_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_296_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_296_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_296_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_297_clock; // @[pe.scala 187:13]
  wire  PE_297_reset; // @[pe.scala 187:13]
  wire  PE_297_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_297_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_297_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_297_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_297_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_297_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_297_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_297_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_297_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_297_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_297_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_298_clock; // @[pe.scala 187:13]
  wire  PE_298_reset; // @[pe.scala 187:13]
  wire  PE_298_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_298_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_298_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_298_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_298_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_298_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_298_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_298_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_298_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_298_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_298_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_299_clock; // @[pe.scala 187:13]
  wire  PE_299_reset; // @[pe.scala 187:13]
  wire  PE_299_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_299_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_299_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_299_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_299_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_299_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_299_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_299_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_299_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_299_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_299_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_300_clock; // @[pe.scala 187:13]
  wire  PE_300_reset; // @[pe.scala 187:13]
  wire  PE_300_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_300_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_300_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_300_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_300_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_300_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_300_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_300_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_300_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_300_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_300_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_301_clock; // @[pe.scala 187:13]
  wire  PE_301_reset; // @[pe.scala 187:13]
  wire  PE_301_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_301_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_301_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_301_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_301_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_301_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_301_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_301_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_301_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_301_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_301_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_302_clock; // @[pe.scala 187:13]
  wire  PE_302_reset; // @[pe.scala 187:13]
  wire  PE_302_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_302_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_302_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_302_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_302_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_302_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_302_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_302_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_302_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_302_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_302_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_303_clock; // @[pe.scala 187:13]
  wire  PE_303_reset; // @[pe.scala 187:13]
  wire  PE_303_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_303_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_303_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_303_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_303_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_303_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_303_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_303_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_303_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_303_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_303_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_304_clock; // @[pe.scala 187:13]
  wire  PE_304_reset; // @[pe.scala 187:13]
  wire  PE_304_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_304_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_304_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_304_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_304_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_304_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_304_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_304_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_304_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_304_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_304_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_305_clock; // @[pe.scala 187:13]
  wire  PE_305_reset; // @[pe.scala 187:13]
  wire  PE_305_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_305_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_305_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_305_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_305_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_305_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_305_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_305_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_305_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_305_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_305_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_306_clock; // @[pe.scala 187:13]
  wire  PE_306_reset; // @[pe.scala 187:13]
  wire  PE_306_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_306_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_306_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_306_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_306_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_306_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_306_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_306_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_306_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_306_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_306_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_307_clock; // @[pe.scala 187:13]
  wire  PE_307_reset; // @[pe.scala 187:13]
  wire  PE_307_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_307_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_307_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_307_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_307_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_307_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_307_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_307_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_307_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_307_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_307_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_308_clock; // @[pe.scala 187:13]
  wire  PE_308_reset; // @[pe.scala 187:13]
  wire  PE_308_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_308_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_308_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_308_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_308_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_308_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_308_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_308_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_308_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_308_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_308_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_309_clock; // @[pe.scala 187:13]
  wire  PE_309_reset; // @[pe.scala 187:13]
  wire  PE_309_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_309_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_309_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_309_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_309_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_309_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_309_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_309_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_309_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_309_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_309_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_310_clock; // @[pe.scala 187:13]
  wire  PE_310_reset; // @[pe.scala 187:13]
  wire  PE_310_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_310_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_310_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_310_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_310_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_310_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_310_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_310_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_310_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_310_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_310_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_311_clock; // @[pe.scala 187:13]
  wire  PE_311_reset; // @[pe.scala 187:13]
  wire  PE_311_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_311_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_311_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_311_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_311_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_311_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_311_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_311_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_311_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_311_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_311_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_312_clock; // @[pe.scala 187:13]
  wire  PE_312_reset; // @[pe.scala 187:13]
  wire  PE_312_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_312_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_312_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_312_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_312_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_312_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_312_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_312_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_312_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_312_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_312_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_313_clock; // @[pe.scala 187:13]
  wire  PE_313_reset; // @[pe.scala 187:13]
  wire  PE_313_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_313_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_313_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_313_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_313_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_313_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_313_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_313_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_313_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_313_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_313_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_314_clock; // @[pe.scala 187:13]
  wire  PE_314_reset; // @[pe.scala 187:13]
  wire  PE_314_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_314_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_314_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_314_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_314_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_314_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_314_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_314_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_314_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_314_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_314_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_315_clock; // @[pe.scala 187:13]
  wire  PE_315_reset; // @[pe.scala 187:13]
  wire  PE_315_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_315_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_315_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_315_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_315_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_315_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_315_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_315_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_315_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_315_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_315_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_316_clock; // @[pe.scala 187:13]
  wire  PE_316_reset; // @[pe.scala 187:13]
  wire  PE_316_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_316_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_316_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_316_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_316_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_316_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_316_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_316_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_316_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_316_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_316_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_317_clock; // @[pe.scala 187:13]
  wire  PE_317_reset; // @[pe.scala 187:13]
  wire  PE_317_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_317_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_317_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_317_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_317_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_317_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_317_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_317_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_317_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_317_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_317_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_318_clock; // @[pe.scala 187:13]
  wire  PE_318_reset; // @[pe.scala 187:13]
  wire  PE_318_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_318_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_318_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_318_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_318_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_318_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_318_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_318_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_318_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_318_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_318_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_319_clock; // @[pe.scala 187:13]
  wire  PE_319_reset; // @[pe.scala 187:13]
  wire  PE_319_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_319_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_319_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_319_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_319_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_319_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_319_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_319_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_319_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_319_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_319_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_320_clock; // @[pe.scala 187:13]
  wire  PE_320_reset; // @[pe.scala 187:13]
  wire  PE_320_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_320_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_320_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_320_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_320_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_320_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_320_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_320_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_320_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_320_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_320_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_321_clock; // @[pe.scala 187:13]
  wire  PE_321_reset; // @[pe.scala 187:13]
  wire  PE_321_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_321_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_321_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_321_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_321_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_321_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_321_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_321_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_321_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_321_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_321_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_322_clock; // @[pe.scala 187:13]
  wire  PE_322_reset; // @[pe.scala 187:13]
  wire  PE_322_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_322_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_322_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_322_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_322_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_322_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_322_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_322_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_322_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_322_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_322_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_323_clock; // @[pe.scala 187:13]
  wire  PE_323_reset; // @[pe.scala 187:13]
  wire  PE_323_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_323_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_323_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_323_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_323_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_323_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_323_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_323_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_323_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_323_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_323_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_324_clock; // @[pe.scala 187:13]
  wire  PE_324_reset; // @[pe.scala 187:13]
  wire  PE_324_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_324_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_324_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_324_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_324_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_324_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_324_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_324_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_324_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_324_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_324_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_325_clock; // @[pe.scala 187:13]
  wire  PE_325_reset; // @[pe.scala 187:13]
  wire  PE_325_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_325_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_325_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_325_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_325_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_325_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_325_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_325_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_325_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_325_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_325_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_326_clock; // @[pe.scala 187:13]
  wire  PE_326_reset; // @[pe.scala 187:13]
  wire  PE_326_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_326_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_326_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_326_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_326_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_326_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_326_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_326_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_326_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_326_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_326_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_327_clock; // @[pe.scala 187:13]
  wire  PE_327_reset; // @[pe.scala 187:13]
  wire  PE_327_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_327_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_327_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_327_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_327_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_327_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_327_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_327_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_327_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_327_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_327_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_328_clock; // @[pe.scala 187:13]
  wire  PE_328_reset; // @[pe.scala 187:13]
  wire  PE_328_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_328_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_328_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_328_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_328_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_328_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_328_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_328_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_328_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_328_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_328_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_329_clock; // @[pe.scala 187:13]
  wire  PE_329_reset; // @[pe.scala 187:13]
  wire  PE_329_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_329_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_329_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_329_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_329_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_329_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_329_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_329_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_329_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_329_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_329_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_330_clock; // @[pe.scala 187:13]
  wire  PE_330_reset; // @[pe.scala 187:13]
  wire  PE_330_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_330_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_330_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_330_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_330_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_330_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_330_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_330_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_330_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_330_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_330_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_331_clock; // @[pe.scala 187:13]
  wire  PE_331_reset; // @[pe.scala 187:13]
  wire  PE_331_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_331_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_331_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_331_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_331_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_331_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_331_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_331_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_331_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_331_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_331_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_332_clock; // @[pe.scala 187:13]
  wire  PE_332_reset; // @[pe.scala 187:13]
  wire  PE_332_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_332_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_332_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_332_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_332_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_332_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_332_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_332_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_332_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_332_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_332_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_333_clock; // @[pe.scala 187:13]
  wire  PE_333_reset; // @[pe.scala 187:13]
  wire  PE_333_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_333_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_333_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_333_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_333_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_333_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_333_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_333_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_333_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_333_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_333_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_334_clock; // @[pe.scala 187:13]
  wire  PE_334_reset; // @[pe.scala 187:13]
  wire  PE_334_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_334_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_334_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_334_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_334_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_334_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_334_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_334_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_334_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_334_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_334_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_335_clock; // @[pe.scala 187:13]
  wire  PE_335_reset; // @[pe.scala 187:13]
  wire  PE_335_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_335_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_335_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_335_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_335_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_335_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_335_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_335_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_335_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_335_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_335_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_336_clock; // @[pe.scala 187:13]
  wire  PE_336_reset; // @[pe.scala 187:13]
  wire  PE_336_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_336_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_336_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_336_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_336_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_336_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_336_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_336_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_336_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_336_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_336_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_337_clock; // @[pe.scala 187:13]
  wire  PE_337_reset; // @[pe.scala 187:13]
  wire  PE_337_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_337_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_337_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_337_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_337_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_337_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_337_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_337_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_337_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_337_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_337_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_338_clock; // @[pe.scala 187:13]
  wire  PE_338_reset; // @[pe.scala 187:13]
  wire  PE_338_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_338_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_338_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_338_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_338_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_338_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_338_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_338_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_338_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_338_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_338_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_339_clock; // @[pe.scala 187:13]
  wire  PE_339_reset; // @[pe.scala 187:13]
  wire  PE_339_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_339_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_339_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_339_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_339_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_339_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_339_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_339_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_339_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_339_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_339_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_340_clock; // @[pe.scala 187:13]
  wire  PE_340_reset; // @[pe.scala 187:13]
  wire  PE_340_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_340_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_340_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_340_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_340_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_340_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_340_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_340_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_340_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_340_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_340_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_341_clock; // @[pe.scala 187:13]
  wire  PE_341_reset; // @[pe.scala 187:13]
  wire  PE_341_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_341_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_341_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_341_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_341_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_341_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_341_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_341_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_341_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_341_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_341_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_342_clock; // @[pe.scala 187:13]
  wire  PE_342_reset; // @[pe.scala 187:13]
  wire  PE_342_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_342_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_342_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_342_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_342_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_342_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_342_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_342_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_342_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_342_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_342_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_343_clock; // @[pe.scala 187:13]
  wire  PE_343_reset; // @[pe.scala 187:13]
  wire  PE_343_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_343_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_343_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_343_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_343_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_343_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_343_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_343_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_343_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_343_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_343_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_344_clock; // @[pe.scala 187:13]
  wire  PE_344_reset; // @[pe.scala 187:13]
  wire  PE_344_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_344_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_344_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_344_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_344_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_344_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_344_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_344_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_344_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_344_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_344_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_345_clock; // @[pe.scala 187:13]
  wire  PE_345_reset; // @[pe.scala 187:13]
  wire  PE_345_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_345_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_345_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_345_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_345_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_345_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_345_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_345_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_345_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_345_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_345_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_346_clock; // @[pe.scala 187:13]
  wire  PE_346_reset; // @[pe.scala 187:13]
  wire  PE_346_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_346_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_346_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_346_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_346_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_346_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_346_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_346_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_346_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_346_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_346_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_347_clock; // @[pe.scala 187:13]
  wire  PE_347_reset; // @[pe.scala 187:13]
  wire  PE_347_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_347_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_347_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_347_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_347_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_347_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_347_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_347_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_347_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_347_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_347_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_348_clock; // @[pe.scala 187:13]
  wire  PE_348_reset; // @[pe.scala 187:13]
  wire  PE_348_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_348_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_348_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_348_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_348_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_348_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_348_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_348_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_348_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_348_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_348_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_349_clock; // @[pe.scala 187:13]
  wire  PE_349_reset; // @[pe.scala 187:13]
  wire  PE_349_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_349_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_349_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_349_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_349_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_349_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_349_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_349_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_349_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_349_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_349_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_350_clock; // @[pe.scala 187:13]
  wire  PE_350_reset; // @[pe.scala 187:13]
  wire  PE_350_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_350_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_350_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_350_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_350_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_350_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_350_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_350_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_350_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_350_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_350_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_351_clock; // @[pe.scala 187:13]
  wire  PE_351_reset; // @[pe.scala 187:13]
  wire  PE_351_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_351_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_351_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_351_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_351_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_351_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_351_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_351_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_351_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_351_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_351_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_352_clock; // @[pe.scala 187:13]
  wire  PE_352_reset; // @[pe.scala 187:13]
  wire  PE_352_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_352_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_352_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_352_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_352_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_352_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_352_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_352_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_352_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_352_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_352_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_353_clock; // @[pe.scala 187:13]
  wire  PE_353_reset; // @[pe.scala 187:13]
  wire  PE_353_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_353_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_353_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_353_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_353_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_353_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_353_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_353_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_353_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_353_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_353_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_354_clock; // @[pe.scala 187:13]
  wire  PE_354_reset; // @[pe.scala 187:13]
  wire  PE_354_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_354_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_354_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_354_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_354_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_354_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_354_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_354_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_354_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_354_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_354_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_355_clock; // @[pe.scala 187:13]
  wire  PE_355_reset; // @[pe.scala 187:13]
  wire  PE_355_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_355_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_355_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_355_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_355_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_355_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_355_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_355_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_355_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_355_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_355_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_356_clock; // @[pe.scala 187:13]
  wire  PE_356_reset; // @[pe.scala 187:13]
  wire  PE_356_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_356_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_356_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_356_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_356_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_356_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_356_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_356_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_356_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_356_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_356_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_357_clock; // @[pe.scala 187:13]
  wire  PE_357_reset; // @[pe.scala 187:13]
  wire  PE_357_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_357_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_357_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_357_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_357_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_357_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_357_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_357_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_357_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_357_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_357_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_358_clock; // @[pe.scala 187:13]
  wire  PE_358_reset; // @[pe.scala 187:13]
  wire  PE_358_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_358_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_358_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_358_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_358_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_358_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_358_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_358_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_358_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_358_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_358_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_359_clock; // @[pe.scala 187:13]
  wire  PE_359_reset; // @[pe.scala 187:13]
  wire  PE_359_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_359_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_359_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_359_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_359_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_359_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_359_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_359_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_359_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_359_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_359_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_360_clock; // @[pe.scala 187:13]
  wire  PE_360_reset; // @[pe.scala 187:13]
  wire  PE_360_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_360_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_360_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_360_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_360_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_360_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_360_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_360_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_360_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_360_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_360_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_361_clock; // @[pe.scala 187:13]
  wire  PE_361_reset; // @[pe.scala 187:13]
  wire  PE_361_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_361_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_361_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_361_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_361_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_361_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_361_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_361_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_361_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_361_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_361_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_362_clock; // @[pe.scala 187:13]
  wire  PE_362_reset; // @[pe.scala 187:13]
  wire  PE_362_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_362_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_362_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_362_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_362_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_362_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_362_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_362_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_362_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_362_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_362_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_363_clock; // @[pe.scala 187:13]
  wire  PE_363_reset; // @[pe.scala 187:13]
  wire  PE_363_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_363_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_363_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_363_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_363_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_363_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_363_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_363_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_363_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_363_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_363_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_364_clock; // @[pe.scala 187:13]
  wire  PE_364_reset; // @[pe.scala 187:13]
  wire  PE_364_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_364_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_364_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_364_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_364_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_364_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_364_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_364_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_364_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_364_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_364_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_365_clock; // @[pe.scala 187:13]
  wire  PE_365_reset; // @[pe.scala 187:13]
  wire  PE_365_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_365_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_365_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_365_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_365_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_365_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_365_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_365_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_365_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_365_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_365_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_366_clock; // @[pe.scala 187:13]
  wire  PE_366_reset; // @[pe.scala 187:13]
  wire  PE_366_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_366_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_366_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_366_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_366_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_366_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_366_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_366_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_366_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_366_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_366_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_367_clock; // @[pe.scala 187:13]
  wire  PE_367_reset; // @[pe.scala 187:13]
  wire  PE_367_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_367_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_367_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_367_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_367_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_367_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_367_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_367_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_367_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_367_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_367_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_368_clock; // @[pe.scala 187:13]
  wire  PE_368_reset; // @[pe.scala 187:13]
  wire  PE_368_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_368_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_368_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_368_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_368_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_368_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_368_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_368_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_368_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_368_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_368_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_369_clock; // @[pe.scala 187:13]
  wire  PE_369_reset; // @[pe.scala 187:13]
  wire  PE_369_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_369_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_369_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_369_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_369_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_369_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_369_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_369_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_369_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_369_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_369_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_370_clock; // @[pe.scala 187:13]
  wire  PE_370_reset; // @[pe.scala 187:13]
  wire  PE_370_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_370_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_370_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_370_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_370_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_370_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_370_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_370_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_370_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_370_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_370_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_371_clock; // @[pe.scala 187:13]
  wire  PE_371_reset; // @[pe.scala 187:13]
  wire  PE_371_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_371_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_371_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_371_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_371_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_371_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_371_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_371_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_371_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_371_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_371_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_372_clock; // @[pe.scala 187:13]
  wire  PE_372_reset; // @[pe.scala 187:13]
  wire  PE_372_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_372_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_372_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_372_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_372_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_372_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_372_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_372_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_372_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_372_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_372_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_373_clock; // @[pe.scala 187:13]
  wire  PE_373_reset; // @[pe.scala 187:13]
  wire  PE_373_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_373_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_373_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_373_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_373_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_373_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_373_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_373_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_373_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_373_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_373_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_374_clock; // @[pe.scala 187:13]
  wire  PE_374_reset; // @[pe.scala 187:13]
  wire  PE_374_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_374_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_374_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_374_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_374_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_374_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_374_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_374_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_374_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_374_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_374_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_375_clock; // @[pe.scala 187:13]
  wire  PE_375_reset; // @[pe.scala 187:13]
  wire  PE_375_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_375_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_375_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_375_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_375_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_375_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_375_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_375_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_375_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_375_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_375_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_376_clock; // @[pe.scala 187:13]
  wire  PE_376_reset; // @[pe.scala 187:13]
  wire  PE_376_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_376_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_376_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_376_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_376_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_376_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_376_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_376_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_376_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_376_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_376_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_377_clock; // @[pe.scala 187:13]
  wire  PE_377_reset; // @[pe.scala 187:13]
  wire  PE_377_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_377_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_377_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_377_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_377_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_377_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_377_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_377_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_377_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_377_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_377_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_378_clock; // @[pe.scala 187:13]
  wire  PE_378_reset; // @[pe.scala 187:13]
  wire  PE_378_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_378_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_378_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_378_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_378_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_378_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_378_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_378_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_378_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_378_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_378_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_379_clock; // @[pe.scala 187:13]
  wire  PE_379_reset; // @[pe.scala 187:13]
  wire  PE_379_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_379_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_379_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_379_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_379_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_379_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_379_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_379_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_379_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_379_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_379_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_380_clock; // @[pe.scala 187:13]
  wire  PE_380_reset; // @[pe.scala 187:13]
  wire  PE_380_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_380_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_380_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_380_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_380_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_380_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_380_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_380_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_380_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_380_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_380_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_381_clock; // @[pe.scala 187:13]
  wire  PE_381_reset; // @[pe.scala 187:13]
  wire  PE_381_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_381_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_381_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_381_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_381_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_381_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_381_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_381_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_381_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_381_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_381_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_382_clock; // @[pe.scala 187:13]
  wire  PE_382_reset; // @[pe.scala 187:13]
  wire  PE_382_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_382_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_382_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_382_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_382_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_382_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_382_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_382_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_382_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_382_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_382_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_383_clock; // @[pe.scala 187:13]
  wire  PE_383_reset; // @[pe.scala 187:13]
  wire  PE_383_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_383_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_383_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_383_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_383_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_383_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_383_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_383_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_383_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_383_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_383_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_384_clock; // @[pe.scala 187:13]
  wire  PE_384_reset; // @[pe.scala 187:13]
  wire  PE_384_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_384_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_384_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_384_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_384_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_384_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_384_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_384_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_384_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_384_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_384_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_385_clock; // @[pe.scala 187:13]
  wire  PE_385_reset; // @[pe.scala 187:13]
  wire  PE_385_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_385_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_385_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_385_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_385_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_385_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_385_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_385_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_385_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_385_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_385_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_386_clock; // @[pe.scala 187:13]
  wire  PE_386_reset; // @[pe.scala 187:13]
  wire  PE_386_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_386_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_386_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_386_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_386_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_386_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_386_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_386_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_386_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_386_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_386_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_387_clock; // @[pe.scala 187:13]
  wire  PE_387_reset; // @[pe.scala 187:13]
  wire  PE_387_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_387_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_387_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_387_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_387_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_387_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_387_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_387_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_387_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_387_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_387_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_388_clock; // @[pe.scala 187:13]
  wire  PE_388_reset; // @[pe.scala 187:13]
  wire  PE_388_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_388_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_388_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_388_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_388_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_388_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_388_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_388_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_388_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_388_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_388_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_389_clock; // @[pe.scala 187:13]
  wire  PE_389_reset; // @[pe.scala 187:13]
  wire  PE_389_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_389_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_389_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_389_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_389_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_389_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_389_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_389_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_389_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_389_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_389_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_390_clock; // @[pe.scala 187:13]
  wire  PE_390_reset; // @[pe.scala 187:13]
  wire  PE_390_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_390_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_390_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_390_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_390_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_390_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_390_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_390_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_390_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_390_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_390_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_391_clock; // @[pe.scala 187:13]
  wire  PE_391_reset; // @[pe.scala 187:13]
  wire  PE_391_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_391_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_391_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_391_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_391_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_391_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_391_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_391_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_391_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_391_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_391_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_392_clock; // @[pe.scala 187:13]
  wire  PE_392_reset; // @[pe.scala 187:13]
  wire  PE_392_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_392_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_392_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_392_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_392_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_392_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_392_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_392_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_392_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_392_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_392_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_393_clock; // @[pe.scala 187:13]
  wire  PE_393_reset; // @[pe.scala 187:13]
  wire  PE_393_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_393_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_393_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_393_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_393_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_393_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_393_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_393_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_393_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_393_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_393_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_394_clock; // @[pe.scala 187:13]
  wire  PE_394_reset; // @[pe.scala 187:13]
  wire  PE_394_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_394_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_394_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_394_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_394_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_394_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_394_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_394_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_394_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_394_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_394_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_395_clock; // @[pe.scala 187:13]
  wire  PE_395_reset; // @[pe.scala 187:13]
  wire  PE_395_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_395_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_395_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_395_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_395_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_395_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_395_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_395_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_395_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_395_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_395_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_396_clock; // @[pe.scala 187:13]
  wire  PE_396_reset; // @[pe.scala 187:13]
  wire  PE_396_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_396_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_396_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_396_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_396_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_396_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_396_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_396_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_396_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_396_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_396_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_397_clock; // @[pe.scala 187:13]
  wire  PE_397_reset; // @[pe.scala 187:13]
  wire  PE_397_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_397_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_397_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_397_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_397_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_397_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_397_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_397_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_397_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_397_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_397_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_398_clock; // @[pe.scala 187:13]
  wire  PE_398_reset; // @[pe.scala 187:13]
  wire  PE_398_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_398_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_398_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_398_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_398_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_398_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_398_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_398_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_398_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_398_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_398_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_399_clock; // @[pe.scala 187:13]
  wire  PE_399_reset; // @[pe.scala 187:13]
  wire  PE_399_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_399_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_399_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_399_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_399_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_399_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_399_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_399_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_399_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_399_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_399_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_400_clock; // @[pe.scala 187:13]
  wire  PE_400_reset; // @[pe.scala 187:13]
  wire  PE_400_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_400_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_400_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_400_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_400_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_400_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_400_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_400_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_400_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_400_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_400_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_401_clock; // @[pe.scala 187:13]
  wire  PE_401_reset; // @[pe.scala 187:13]
  wire  PE_401_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_401_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_401_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_401_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_401_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_401_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_401_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_401_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_401_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_401_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_401_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_402_clock; // @[pe.scala 187:13]
  wire  PE_402_reset; // @[pe.scala 187:13]
  wire  PE_402_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_402_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_402_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_402_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_402_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_402_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_402_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_402_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_402_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_402_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_402_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_403_clock; // @[pe.scala 187:13]
  wire  PE_403_reset; // @[pe.scala 187:13]
  wire  PE_403_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_403_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_403_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_403_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_403_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_403_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_403_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_403_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_403_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_403_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_403_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_404_clock; // @[pe.scala 187:13]
  wire  PE_404_reset; // @[pe.scala 187:13]
  wire  PE_404_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_404_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_404_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_404_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_404_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_404_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_404_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_404_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_404_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_404_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_404_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_405_clock; // @[pe.scala 187:13]
  wire  PE_405_reset; // @[pe.scala 187:13]
  wire  PE_405_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_405_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_405_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_405_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_405_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_405_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_405_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_405_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_405_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_405_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_405_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_406_clock; // @[pe.scala 187:13]
  wire  PE_406_reset; // @[pe.scala 187:13]
  wire  PE_406_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_406_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_406_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_406_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_406_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_406_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_406_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_406_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_406_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_406_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_406_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_407_clock; // @[pe.scala 187:13]
  wire  PE_407_reset; // @[pe.scala 187:13]
  wire  PE_407_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_407_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_407_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_407_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_407_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_407_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_407_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_407_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_407_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_407_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_407_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_408_clock; // @[pe.scala 187:13]
  wire  PE_408_reset; // @[pe.scala 187:13]
  wire  PE_408_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_408_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_408_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_408_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_408_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_408_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_408_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_408_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_408_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_408_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_408_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_409_clock; // @[pe.scala 187:13]
  wire  PE_409_reset; // @[pe.scala 187:13]
  wire  PE_409_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_409_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_409_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_409_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_409_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_409_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_409_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_409_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_409_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_409_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_409_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_410_clock; // @[pe.scala 187:13]
  wire  PE_410_reset; // @[pe.scala 187:13]
  wire  PE_410_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_410_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_410_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_410_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_410_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_410_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_410_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_410_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_410_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_410_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_410_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_411_clock; // @[pe.scala 187:13]
  wire  PE_411_reset; // @[pe.scala 187:13]
  wire  PE_411_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_411_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_411_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_411_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_411_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_411_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_411_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_411_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_411_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_411_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_411_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_412_clock; // @[pe.scala 187:13]
  wire  PE_412_reset; // @[pe.scala 187:13]
  wire  PE_412_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_412_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_412_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_412_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_412_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_412_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_412_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_412_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_412_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_412_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_412_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_413_clock; // @[pe.scala 187:13]
  wire  PE_413_reset; // @[pe.scala 187:13]
  wire  PE_413_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_413_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_413_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_413_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_413_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_413_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_413_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_413_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_413_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_413_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_413_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_414_clock; // @[pe.scala 187:13]
  wire  PE_414_reset; // @[pe.scala 187:13]
  wire  PE_414_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_414_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_414_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_414_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_414_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_414_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_414_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_414_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_414_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_414_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_414_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_415_clock; // @[pe.scala 187:13]
  wire  PE_415_reset; // @[pe.scala 187:13]
  wire  PE_415_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_415_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_415_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_415_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_415_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_415_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_415_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_415_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_415_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_415_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_415_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_416_clock; // @[pe.scala 187:13]
  wire  PE_416_reset; // @[pe.scala 187:13]
  wire  PE_416_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_416_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_416_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_416_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_416_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_416_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_416_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_416_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_416_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_416_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_416_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_417_clock; // @[pe.scala 187:13]
  wire  PE_417_reset; // @[pe.scala 187:13]
  wire  PE_417_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_417_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_417_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_417_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_417_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_417_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_417_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_417_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_417_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_417_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_417_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_418_clock; // @[pe.scala 187:13]
  wire  PE_418_reset; // @[pe.scala 187:13]
  wire  PE_418_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_418_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_418_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_418_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_418_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_418_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_418_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_418_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_418_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_418_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_418_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_419_clock; // @[pe.scala 187:13]
  wire  PE_419_reset; // @[pe.scala 187:13]
  wire  PE_419_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_419_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_419_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_419_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_419_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_419_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_419_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_419_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_419_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_419_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_419_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_420_clock; // @[pe.scala 187:13]
  wire  PE_420_reset; // @[pe.scala 187:13]
  wire  PE_420_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_420_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_420_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_420_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_420_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_420_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_420_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_420_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_420_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_420_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_420_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_421_clock; // @[pe.scala 187:13]
  wire  PE_421_reset; // @[pe.scala 187:13]
  wire  PE_421_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_421_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_421_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_421_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_421_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_421_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_421_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_421_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_421_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_421_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_421_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_422_clock; // @[pe.scala 187:13]
  wire  PE_422_reset; // @[pe.scala 187:13]
  wire  PE_422_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_422_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_422_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_422_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_422_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_422_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_422_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_422_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_422_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_422_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_422_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_423_clock; // @[pe.scala 187:13]
  wire  PE_423_reset; // @[pe.scala 187:13]
  wire  PE_423_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_423_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_423_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_423_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_423_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_423_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_423_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_423_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_423_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_423_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_423_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_424_clock; // @[pe.scala 187:13]
  wire  PE_424_reset; // @[pe.scala 187:13]
  wire  PE_424_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_424_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_424_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_424_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_424_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_424_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_424_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_424_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_424_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_424_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_424_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_425_clock; // @[pe.scala 187:13]
  wire  PE_425_reset; // @[pe.scala 187:13]
  wire  PE_425_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_425_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_425_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_425_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_425_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_425_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_425_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_425_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_425_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_425_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_425_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_426_clock; // @[pe.scala 187:13]
  wire  PE_426_reset; // @[pe.scala 187:13]
  wire  PE_426_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_426_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_426_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_426_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_426_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_426_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_426_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_426_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_426_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_426_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_426_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_427_clock; // @[pe.scala 187:13]
  wire  PE_427_reset; // @[pe.scala 187:13]
  wire  PE_427_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_427_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_427_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_427_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_427_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_427_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_427_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_427_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_427_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_427_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_427_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_428_clock; // @[pe.scala 187:13]
  wire  PE_428_reset; // @[pe.scala 187:13]
  wire  PE_428_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_428_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_428_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_428_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_428_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_428_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_428_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_428_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_428_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_428_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_428_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_429_clock; // @[pe.scala 187:13]
  wire  PE_429_reset; // @[pe.scala 187:13]
  wire  PE_429_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_429_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_429_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_429_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_429_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_429_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_429_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_429_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_429_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_429_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_429_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_430_clock; // @[pe.scala 187:13]
  wire  PE_430_reset; // @[pe.scala 187:13]
  wire  PE_430_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_430_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_430_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_430_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_430_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_430_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_430_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_430_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_430_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_430_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_430_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_431_clock; // @[pe.scala 187:13]
  wire  PE_431_reset; // @[pe.scala 187:13]
  wire  PE_431_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_431_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_431_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_431_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_431_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_431_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_431_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_431_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_431_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_431_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_431_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_432_clock; // @[pe.scala 187:13]
  wire  PE_432_reset; // @[pe.scala 187:13]
  wire  PE_432_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_432_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_432_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_432_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_432_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_432_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_432_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_432_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_432_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_432_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_432_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_433_clock; // @[pe.scala 187:13]
  wire  PE_433_reset; // @[pe.scala 187:13]
  wire  PE_433_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_433_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_433_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_433_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_433_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_433_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_433_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_433_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_433_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_433_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_433_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_434_clock; // @[pe.scala 187:13]
  wire  PE_434_reset; // @[pe.scala 187:13]
  wire  PE_434_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_434_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_434_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_434_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_434_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_434_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_434_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_434_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_434_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_434_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_434_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_435_clock; // @[pe.scala 187:13]
  wire  PE_435_reset; // @[pe.scala 187:13]
  wire  PE_435_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_435_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_435_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_435_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_435_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_435_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_435_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_435_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_435_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_435_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_435_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_436_clock; // @[pe.scala 187:13]
  wire  PE_436_reset; // @[pe.scala 187:13]
  wire  PE_436_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_436_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_436_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_436_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_436_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_436_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_436_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_436_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_436_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_436_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_436_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_437_clock; // @[pe.scala 187:13]
  wire  PE_437_reset; // @[pe.scala 187:13]
  wire  PE_437_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_437_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_437_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_437_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_437_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_437_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_437_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_437_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_437_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_437_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_437_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_438_clock; // @[pe.scala 187:13]
  wire  PE_438_reset; // @[pe.scala 187:13]
  wire  PE_438_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_438_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_438_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_438_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_438_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_438_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_438_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_438_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_438_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_438_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_438_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_439_clock; // @[pe.scala 187:13]
  wire  PE_439_reset; // @[pe.scala 187:13]
  wire  PE_439_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_439_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_439_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_439_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_439_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_439_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_439_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_439_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_439_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_439_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_439_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_440_clock; // @[pe.scala 187:13]
  wire  PE_440_reset; // @[pe.scala 187:13]
  wire  PE_440_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_440_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_440_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_440_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_440_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_440_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_440_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_440_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_440_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_440_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_440_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_441_clock; // @[pe.scala 187:13]
  wire  PE_441_reset; // @[pe.scala 187:13]
  wire  PE_441_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_441_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_441_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_441_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_441_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_441_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_441_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_441_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_441_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_441_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_441_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_442_clock; // @[pe.scala 187:13]
  wire  PE_442_reset; // @[pe.scala 187:13]
  wire  PE_442_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_442_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_442_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_442_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_442_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_442_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_442_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_442_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_442_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_442_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_442_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_443_clock; // @[pe.scala 187:13]
  wire  PE_443_reset; // @[pe.scala 187:13]
  wire  PE_443_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_443_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_443_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_443_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_443_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_443_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_443_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_443_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_443_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_443_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_443_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_444_clock; // @[pe.scala 187:13]
  wire  PE_444_reset; // @[pe.scala 187:13]
  wire  PE_444_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_444_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_444_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_444_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_444_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_444_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_444_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_444_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_444_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_444_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_444_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_445_clock; // @[pe.scala 187:13]
  wire  PE_445_reset; // @[pe.scala 187:13]
  wire  PE_445_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_445_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_445_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_445_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_445_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_445_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_445_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_445_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_445_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_445_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_445_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_446_clock; // @[pe.scala 187:13]
  wire  PE_446_reset; // @[pe.scala 187:13]
  wire  PE_446_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_446_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_446_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_446_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_446_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_446_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_446_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_446_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_446_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_446_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_446_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_447_clock; // @[pe.scala 187:13]
  wire  PE_447_reset; // @[pe.scala 187:13]
  wire  PE_447_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_447_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_447_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_447_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_447_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_447_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_447_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_447_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_447_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_447_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_447_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_448_clock; // @[pe.scala 187:13]
  wire  PE_448_reset; // @[pe.scala 187:13]
  wire  PE_448_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_448_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_448_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_448_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_448_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_448_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_448_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_448_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_448_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_448_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_448_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_449_clock; // @[pe.scala 187:13]
  wire  PE_449_reset; // @[pe.scala 187:13]
  wire  PE_449_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_449_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_449_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_449_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_449_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_449_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_449_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_449_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_449_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_449_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_449_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_450_clock; // @[pe.scala 187:13]
  wire  PE_450_reset; // @[pe.scala 187:13]
  wire  PE_450_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_450_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_450_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_450_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_450_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_450_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_450_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_450_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_450_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_450_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_450_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_451_clock; // @[pe.scala 187:13]
  wire  PE_451_reset; // @[pe.scala 187:13]
  wire  PE_451_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_451_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_451_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_451_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_451_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_451_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_451_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_451_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_451_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_451_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_451_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_452_clock; // @[pe.scala 187:13]
  wire  PE_452_reset; // @[pe.scala 187:13]
  wire  PE_452_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_452_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_452_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_452_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_452_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_452_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_452_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_452_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_452_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_452_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_452_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_453_clock; // @[pe.scala 187:13]
  wire  PE_453_reset; // @[pe.scala 187:13]
  wire  PE_453_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_453_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_453_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_453_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_453_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_453_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_453_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_453_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_453_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_453_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_453_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_454_clock; // @[pe.scala 187:13]
  wire  PE_454_reset; // @[pe.scala 187:13]
  wire  PE_454_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_454_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_454_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_454_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_454_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_454_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_454_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_454_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_454_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_454_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_454_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_455_clock; // @[pe.scala 187:13]
  wire  PE_455_reset; // @[pe.scala 187:13]
  wire  PE_455_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_455_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_455_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_455_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_455_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_455_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_455_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_455_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_455_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_455_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_455_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_456_clock; // @[pe.scala 187:13]
  wire  PE_456_reset; // @[pe.scala 187:13]
  wire  PE_456_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_456_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_456_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_456_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_456_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_456_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_456_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_456_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_456_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_456_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_456_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_457_clock; // @[pe.scala 187:13]
  wire  PE_457_reset; // @[pe.scala 187:13]
  wire  PE_457_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_457_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_457_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_457_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_457_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_457_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_457_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_457_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_457_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_457_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_457_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_458_clock; // @[pe.scala 187:13]
  wire  PE_458_reset; // @[pe.scala 187:13]
  wire  PE_458_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_458_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_458_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_458_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_458_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_458_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_458_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_458_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_458_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_458_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_458_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_459_clock; // @[pe.scala 187:13]
  wire  PE_459_reset; // @[pe.scala 187:13]
  wire  PE_459_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_459_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_459_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_459_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_459_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_459_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_459_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_459_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_459_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_459_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_459_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_460_clock; // @[pe.scala 187:13]
  wire  PE_460_reset; // @[pe.scala 187:13]
  wire  PE_460_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_460_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_460_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_460_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_460_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_460_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_460_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_460_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_460_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_460_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_460_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_461_clock; // @[pe.scala 187:13]
  wire  PE_461_reset; // @[pe.scala 187:13]
  wire  PE_461_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_461_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_461_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_461_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_461_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_461_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_461_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_461_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_461_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_461_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_461_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_462_clock; // @[pe.scala 187:13]
  wire  PE_462_reset; // @[pe.scala 187:13]
  wire  PE_462_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_462_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_462_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_462_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_462_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_462_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_462_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_462_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_462_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_462_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_462_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_463_clock; // @[pe.scala 187:13]
  wire  PE_463_reset; // @[pe.scala 187:13]
  wire  PE_463_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_463_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_463_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_463_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_463_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_463_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_463_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_463_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_463_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_463_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_463_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_464_clock; // @[pe.scala 187:13]
  wire  PE_464_reset; // @[pe.scala 187:13]
  wire  PE_464_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_464_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_464_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_464_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_464_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_464_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_464_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_464_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_464_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_464_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_464_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_465_clock; // @[pe.scala 187:13]
  wire  PE_465_reset; // @[pe.scala 187:13]
  wire  PE_465_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_465_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_465_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_465_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_465_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_465_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_465_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_465_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_465_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_465_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_465_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_466_clock; // @[pe.scala 187:13]
  wire  PE_466_reset; // @[pe.scala 187:13]
  wire  PE_466_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_466_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_466_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_466_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_466_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_466_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_466_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_466_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_466_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_466_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_466_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_467_clock; // @[pe.scala 187:13]
  wire  PE_467_reset; // @[pe.scala 187:13]
  wire  PE_467_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_467_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_467_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_467_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_467_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_467_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_467_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_467_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_467_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_467_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_467_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_468_clock; // @[pe.scala 187:13]
  wire  PE_468_reset; // @[pe.scala 187:13]
  wire  PE_468_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_468_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_468_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_468_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_468_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_468_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_468_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_468_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_468_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_468_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_468_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_469_clock; // @[pe.scala 187:13]
  wire  PE_469_reset; // @[pe.scala 187:13]
  wire  PE_469_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_469_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_469_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_469_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_469_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_469_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_469_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_469_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_469_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_469_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_469_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_470_clock; // @[pe.scala 187:13]
  wire  PE_470_reset; // @[pe.scala 187:13]
  wire  PE_470_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_470_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_470_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_470_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_470_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_470_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_470_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_470_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_470_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_470_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_470_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_471_clock; // @[pe.scala 187:13]
  wire  PE_471_reset; // @[pe.scala 187:13]
  wire  PE_471_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_471_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_471_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_471_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_471_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_471_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_471_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_471_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_471_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_471_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_471_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_472_clock; // @[pe.scala 187:13]
  wire  PE_472_reset; // @[pe.scala 187:13]
  wire  PE_472_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_472_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_472_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_472_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_472_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_472_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_472_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_472_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_472_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_472_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_472_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_473_clock; // @[pe.scala 187:13]
  wire  PE_473_reset; // @[pe.scala 187:13]
  wire  PE_473_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_473_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_473_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_473_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_473_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_473_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_473_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_473_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_473_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_473_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_473_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_474_clock; // @[pe.scala 187:13]
  wire  PE_474_reset; // @[pe.scala 187:13]
  wire  PE_474_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_474_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_474_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_474_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_474_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_474_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_474_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_474_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_474_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_474_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_474_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_475_clock; // @[pe.scala 187:13]
  wire  PE_475_reset; // @[pe.scala 187:13]
  wire  PE_475_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_475_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_475_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_475_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_475_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_475_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_475_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_475_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_475_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_475_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_475_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_476_clock; // @[pe.scala 187:13]
  wire  PE_476_reset; // @[pe.scala 187:13]
  wire  PE_476_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_476_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_476_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_476_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_476_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_476_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_476_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_476_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_476_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_476_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_476_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_477_clock; // @[pe.scala 187:13]
  wire  PE_477_reset; // @[pe.scala 187:13]
  wire  PE_477_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_477_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_477_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_477_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_477_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_477_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_477_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_477_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_477_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_477_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_477_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_478_clock; // @[pe.scala 187:13]
  wire  PE_478_reset; // @[pe.scala 187:13]
  wire  PE_478_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_478_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_478_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_478_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_478_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_478_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_478_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_478_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_478_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_478_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_478_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_479_clock; // @[pe.scala 187:13]
  wire  PE_479_reset; // @[pe.scala 187:13]
  wire  PE_479_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_479_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_479_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_479_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_479_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_479_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_479_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_479_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_479_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_479_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_479_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_480_clock; // @[pe.scala 187:13]
  wire  PE_480_reset; // @[pe.scala 187:13]
  wire  PE_480_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_480_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_480_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_480_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_480_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_480_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_480_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_480_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_480_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_480_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_480_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_481_clock; // @[pe.scala 187:13]
  wire  PE_481_reset; // @[pe.scala 187:13]
  wire  PE_481_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_481_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_481_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_481_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_481_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_481_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_481_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_481_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_481_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_481_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_481_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_482_clock; // @[pe.scala 187:13]
  wire  PE_482_reset; // @[pe.scala 187:13]
  wire  PE_482_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_482_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_482_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_482_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_482_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_482_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_482_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_482_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_482_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_482_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_482_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_483_clock; // @[pe.scala 187:13]
  wire  PE_483_reset; // @[pe.scala 187:13]
  wire  PE_483_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_483_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_483_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_483_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_483_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_483_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_483_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_483_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_483_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_483_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_483_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_484_clock; // @[pe.scala 187:13]
  wire  PE_484_reset; // @[pe.scala 187:13]
  wire  PE_484_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_484_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_484_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_484_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_484_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_484_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_484_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_484_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_484_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_484_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_484_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_485_clock; // @[pe.scala 187:13]
  wire  PE_485_reset; // @[pe.scala 187:13]
  wire  PE_485_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_485_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_485_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_485_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_485_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_485_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_485_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_485_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_485_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_485_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_485_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_486_clock; // @[pe.scala 187:13]
  wire  PE_486_reset; // @[pe.scala 187:13]
  wire  PE_486_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_486_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_486_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_486_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_486_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_486_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_486_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_486_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_486_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_486_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_486_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_487_clock; // @[pe.scala 187:13]
  wire  PE_487_reset; // @[pe.scala 187:13]
  wire  PE_487_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_487_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_487_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_487_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_487_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_487_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_487_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_487_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_487_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_487_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_487_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_488_clock; // @[pe.scala 187:13]
  wire  PE_488_reset; // @[pe.scala 187:13]
  wire  PE_488_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_488_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_488_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_488_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_488_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_488_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_488_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_488_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_488_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_488_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_488_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_489_clock; // @[pe.scala 187:13]
  wire  PE_489_reset; // @[pe.scala 187:13]
  wire  PE_489_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_489_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_489_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_489_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_489_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_489_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_489_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_489_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_489_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_489_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_489_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_490_clock; // @[pe.scala 187:13]
  wire  PE_490_reset; // @[pe.scala 187:13]
  wire  PE_490_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_490_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_490_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_490_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_490_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_490_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_490_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_490_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_490_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_490_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_490_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_491_clock; // @[pe.scala 187:13]
  wire  PE_491_reset; // @[pe.scala 187:13]
  wire  PE_491_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_491_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_491_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_491_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_491_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_491_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_491_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_491_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_491_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_491_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_491_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_492_clock; // @[pe.scala 187:13]
  wire  PE_492_reset; // @[pe.scala 187:13]
  wire  PE_492_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_492_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_492_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_492_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_492_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_492_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_492_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_492_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_492_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_492_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_492_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_493_clock; // @[pe.scala 187:13]
  wire  PE_493_reset; // @[pe.scala 187:13]
  wire  PE_493_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_493_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_493_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_493_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_493_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_493_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_493_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_493_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_493_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_493_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_493_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_494_clock; // @[pe.scala 187:13]
  wire  PE_494_reset; // @[pe.scala 187:13]
  wire  PE_494_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_494_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_494_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_494_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_494_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_494_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_494_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_494_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_494_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_494_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_494_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_495_clock; // @[pe.scala 187:13]
  wire  PE_495_reset; // @[pe.scala 187:13]
  wire  PE_495_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_495_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_495_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_495_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_495_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_495_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_495_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_495_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_495_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_495_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_495_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_496_clock; // @[pe.scala 187:13]
  wire  PE_496_reset; // @[pe.scala 187:13]
  wire  PE_496_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_496_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_496_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_496_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_496_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_496_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_496_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_496_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_496_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_496_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_496_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_497_clock; // @[pe.scala 187:13]
  wire  PE_497_reset; // @[pe.scala 187:13]
  wire  PE_497_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_497_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_497_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_497_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_497_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_497_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_497_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_497_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_497_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_497_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_497_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_498_clock; // @[pe.scala 187:13]
  wire  PE_498_reset; // @[pe.scala 187:13]
  wire  PE_498_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_498_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_498_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_498_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_498_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_498_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_498_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_498_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_498_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_498_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_498_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_499_clock; // @[pe.scala 187:13]
  wire  PE_499_reset; // @[pe.scala 187:13]
  wire  PE_499_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_499_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_499_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_499_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_499_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_499_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_499_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_499_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_499_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_499_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_499_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_500_clock; // @[pe.scala 187:13]
  wire  PE_500_reset; // @[pe.scala 187:13]
  wire  PE_500_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_500_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_500_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_500_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_500_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_500_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_500_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_500_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_500_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_500_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_500_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_501_clock; // @[pe.scala 187:13]
  wire  PE_501_reset; // @[pe.scala 187:13]
  wire  PE_501_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_501_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_501_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_501_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_501_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_501_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_501_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_501_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_501_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_501_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_501_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_502_clock; // @[pe.scala 187:13]
  wire  PE_502_reset; // @[pe.scala 187:13]
  wire  PE_502_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_502_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_502_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_502_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_502_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_502_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_502_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_502_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_502_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_502_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_502_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_503_clock; // @[pe.scala 187:13]
  wire  PE_503_reset; // @[pe.scala 187:13]
  wire  PE_503_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_503_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_503_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_503_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_503_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_503_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_503_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_503_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_503_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_503_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_503_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_504_clock; // @[pe.scala 187:13]
  wire  PE_504_reset; // @[pe.scala 187:13]
  wire  PE_504_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_504_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_504_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_504_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_504_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_504_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_504_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_504_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_504_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_504_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_504_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_505_clock; // @[pe.scala 187:13]
  wire  PE_505_reset; // @[pe.scala 187:13]
  wire  PE_505_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_505_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_505_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_505_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_505_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_505_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_505_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_505_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_505_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_505_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_505_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_506_clock; // @[pe.scala 187:13]
  wire  PE_506_reset; // @[pe.scala 187:13]
  wire  PE_506_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_506_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_506_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_506_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_506_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_506_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_506_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_506_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_506_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_506_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_506_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_507_clock; // @[pe.scala 187:13]
  wire  PE_507_reset; // @[pe.scala 187:13]
  wire  PE_507_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_507_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_507_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_507_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_507_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_507_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_507_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_507_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_507_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_507_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_507_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_508_clock; // @[pe.scala 187:13]
  wire  PE_508_reset; // @[pe.scala 187:13]
  wire  PE_508_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_508_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_508_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_508_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_508_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_508_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_508_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_508_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_508_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_508_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_508_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_509_clock; // @[pe.scala 187:13]
  wire  PE_509_reset; // @[pe.scala 187:13]
  wire  PE_509_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_509_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_509_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_509_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_509_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_509_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_509_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_509_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_509_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_509_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_509_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_510_clock; // @[pe.scala 187:13]
  wire  PE_510_reset; // @[pe.scala 187:13]
  wire  PE_510_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_510_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_510_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_510_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_510_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_510_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_510_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_510_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_510_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_510_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_510_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_511_clock; // @[pe.scala 187:13]
  wire  PE_511_reset; // @[pe.scala 187:13]
  wire  PE_511_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_511_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_511_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_511_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_511_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_511_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_511_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_511_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_511_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_511_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_511_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_512_clock; // @[pe.scala 187:13]
  wire  PE_512_reset; // @[pe.scala 187:13]
  wire  PE_512_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_512_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_512_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_512_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_512_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_512_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_512_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_512_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_512_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_512_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_512_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_513_clock; // @[pe.scala 187:13]
  wire  PE_513_reset; // @[pe.scala 187:13]
  wire  PE_513_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_513_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_513_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_513_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_513_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_513_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_513_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_513_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_513_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_513_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_513_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_514_clock; // @[pe.scala 187:13]
  wire  PE_514_reset; // @[pe.scala 187:13]
  wire  PE_514_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_514_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_514_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_514_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_514_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_514_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_514_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_514_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_514_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_514_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_514_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_515_clock; // @[pe.scala 187:13]
  wire  PE_515_reset; // @[pe.scala 187:13]
  wire  PE_515_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_515_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_515_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_515_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_515_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_515_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_515_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_515_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_515_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_515_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_515_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_516_clock; // @[pe.scala 187:13]
  wire  PE_516_reset; // @[pe.scala 187:13]
  wire  PE_516_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_516_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_516_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_516_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_516_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_516_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_516_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_516_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_516_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_516_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_516_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_517_clock; // @[pe.scala 187:13]
  wire  PE_517_reset; // @[pe.scala 187:13]
  wire  PE_517_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_517_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_517_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_517_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_517_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_517_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_517_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_517_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_517_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_517_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_517_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_518_clock; // @[pe.scala 187:13]
  wire  PE_518_reset; // @[pe.scala 187:13]
  wire  PE_518_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_518_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_518_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_518_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_518_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_518_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_518_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_518_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_518_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_518_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_518_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_519_clock; // @[pe.scala 187:13]
  wire  PE_519_reset; // @[pe.scala 187:13]
  wire  PE_519_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_519_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_519_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_519_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_519_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_519_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_519_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_519_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_519_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_519_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_519_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_520_clock; // @[pe.scala 187:13]
  wire  PE_520_reset; // @[pe.scala 187:13]
  wire  PE_520_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_520_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_520_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_520_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_520_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_520_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_520_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_520_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_520_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_520_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_520_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_521_clock; // @[pe.scala 187:13]
  wire  PE_521_reset; // @[pe.scala 187:13]
  wire  PE_521_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_521_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_521_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_521_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_521_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_521_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_521_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_521_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_521_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_521_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_521_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_522_clock; // @[pe.scala 187:13]
  wire  PE_522_reset; // @[pe.scala 187:13]
  wire  PE_522_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_522_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_522_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_522_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_522_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_522_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_522_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_522_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_522_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_522_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_522_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_523_clock; // @[pe.scala 187:13]
  wire  PE_523_reset; // @[pe.scala 187:13]
  wire  PE_523_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_523_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_523_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_523_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_523_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_523_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_523_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_523_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_523_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_523_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_523_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_524_clock; // @[pe.scala 187:13]
  wire  PE_524_reset; // @[pe.scala 187:13]
  wire  PE_524_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_524_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_524_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_524_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_524_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_524_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_524_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_524_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_524_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_524_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_524_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_525_clock; // @[pe.scala 187:13]
  wire  PE_525_reset; // @[pe.scala 187:13]
  wire  PE_525_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_525_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_525_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_525_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_525_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_525_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_525_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_525_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_525_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_525_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_525_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_526_clock; // @[pe.scala 187:13]
  wire  PE_526_reset; // @[pe.scala 187:13]
  wire  PE_526_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_526_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_526_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_526_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_526_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_526_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_526_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_526_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_526_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_526_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_526_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_527_clock; // @[pe.scala 187:13]
  wire  PE_527_reset; // @[pe.scala 187:13]
  wire  PE_527_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_527_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_527_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_527_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_527_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_527_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_527_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_527_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_527_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_527_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_527_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_528_clock; // @[pe.scala 187:13]
  wire  PE_528_reset; // @[pe.scala 187:13]
  wire  PE_528_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_528_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_528_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_528_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_528_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_528_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_528_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_528_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_528_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_528_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_528_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_529_clock; // @[pe.scala 187:13]
  wire  PE_529_reset; // @[pe.scala 187:13]
  wire  PE_529_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_529_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_529_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_529_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_529_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_529_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_529_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_529_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_529_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_529_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_529_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_530_clock; // @[pe.scala 187:13]
  wire  PE_530_reset; // @[pe.scala 187:13]
  wire  PE_530_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_530_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_530_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_530_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_530_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_530_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_530_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_530_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_530_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_530_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_530_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_531_clock; // @[pe.scala 187:13]
  wire  PE_531_reset; // @[pe.scala 187:13]
  wire  PE_531_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_531_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_531_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_531_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_531_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_531_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_531_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_531_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_531_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_531_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_531_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_532_clock; // @[pe.scala 187:13]
  wire  PE_532_reset; // @[pe.scala 187:13]
  wire  PE_532_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_532_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_532_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_532_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_532_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_532_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_532_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_532_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_532_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_532_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_532_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_533_clock; // @[pe.scala 187:13]
  wire  PE_533_reset; // @[pe.scala 187:13]
  wire  PE_533_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_533_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_533_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_533_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_533_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_533_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_533_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_533_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_533_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_533_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_533_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_534_clock; // @[pe.scala 187:13]
  wire  PE_534_reset; // @[pe.scala 187:13]
  wire  PE_534_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_534_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_534_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_534_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_534_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_534_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_534_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_534_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_534_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_534_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_534_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_535_clock; // @[pe.scala 187:13]
  wire  PE_535_reset; // @[pe.scala 187:13]
  wire  PE_535_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_535_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_535_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_535_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_535_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_535_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_535_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_535_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_535_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_535_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_535_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_536_clock; // @[pe.scala 187:13]
  wire  PE_536_reset; // @[pe.scala 187:13]
  wire  PE_536_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_536_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_536_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_536_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_536_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_536_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_536_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_536_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_536_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_536_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_536_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_537_clock; // @[pe.scala 187:13]
  wire  PE_537_reset; // @[pe.scala 187:13]
  wire  PE_537_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_537_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_537_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_537_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_537_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_537_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_537_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_537_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_537_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_537_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_537_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_538_clock; // @[pe.scala 187:13]
  wire  PE_538_reset; // @[pe.scala 187:13]
  wire  PE_538_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_538_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_538_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_538_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_538_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_538_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_538_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_538_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_538_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_538_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_538_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_539_clock; // @[pe.scala 187:13]
  wire  PE_539_reset; // @[pe.scala 187:13]
  wire  PE_539_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_539_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_539_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_539_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_539_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_539_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_539_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_539_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_539_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_539_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_539_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_540_clock; // @[pe.scala 187:13]
  wire  PE_540_reset; // @[pe.scala 187:13]
  wire  PE_540_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_540_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_540_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_540_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_540_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_540_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_540_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_540_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_540_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_540_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_540_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_541_clock; // @[pe.scala 187:13]
  wire  PE_541_reset; // @[pe.scala 187:13]
  wire  PE_541_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_541_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_541_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_541_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_541_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_541_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_541_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_541_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_541_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_541_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_541_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_542_clock; // @[pe.scala 187:13]
  wire  PE_542_reset; // @[pe.scala 187:13]
  wire  PE_542_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_542_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_542_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_542_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_542_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_542_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_542_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_542_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_542_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_542_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_542_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_543_clock; // @[pe.scala 187:13]
  wire  PE_543_reset; // @[pe.scala 187:13]
  wire  PE_543_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_543_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_543_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_543_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_543_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_543_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_543_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_543_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_543_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_543_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_543_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_544_clock; // @[pe.scala 187:13]
  wire  PE_544_reset; // @[pe.scala 187:13]
  wire  PE_544_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_544_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_544_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_544_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_544_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_544_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_544_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_544_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_544_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_544_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_544_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_545_clock; // @[pe.scala 187:13]
  wire  PE_545_reset; // @[pe.scala 187:13]
  wire  PE_545_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_545_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_545_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_545_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_545_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_545_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_545_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_545_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_545_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_545_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_545_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_546_clock; // @[pe.scala 187:13]
  wire  PE_546_reset; // @[pe.scala 187:13]
  wire  PE_546_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_546_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_546_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_546_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_546_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_546_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_546_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_546_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_546_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_546_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_546_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_547_clock; // @[pe.scala 187:13]
  wire  PE_547_reset; // @[pe.scala 187:13]
  wire  PE_547_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_547_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_547_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_547_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_547_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_547_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_547_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_547_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_547_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_547_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_547_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_548_clock; // @[pe.scala 187:13]
  wire  PE_548_reset; // @[pe.scala 187:13]
  wire  PE_548_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_548_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_548_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_548_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_548_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_548_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_548_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_548_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_548_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_548_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_548_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_549_clock; // @[pe.scala 187:13]
  wire  PE_549_reset; // @[pe.scala 187:13]
  wire  PE_549_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_549_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_549_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_549_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_549_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_549_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_549_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_549_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_549_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_549_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_549_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_550_clock; // @[pe.scala 187:13]
  wire  PE_550_reset; // @[pe.scala 187:13]
  wire  PE_550_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_550_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_550_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_550_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_550_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_550_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_550_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_550_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_550_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_550_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_550_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_551_clock; // @[pe.scala 187:13]
  wire  PE_551_reset; // @[pe.scala 187:13]
  wire  PE_551_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_551_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_551_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_551_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_551_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_551_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_551_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_551_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_551_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_551_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_551_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_552_clock; // @[pe.scala 187:13]
  wire  PE_552_reset; // @[pe.scala 187:13]
  wire  PE_552_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_552_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_552_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_552_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_552_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_552_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_552_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_552_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_552_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_552_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_552_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_553_clock; // @[pe.scala 187:13]
  wire  PE_553_reset; // @[pe.scala 187:13]
  wire  PE_553_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_553_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_553_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_553_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_553_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_553_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_553_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_553_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_553_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_553_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_553_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_554_clock; // @[pe.scala 187:13]
  wire  PE_554_reset; // @[pe.scala 187:13]
  wire  PE_554_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_554_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_554_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_554_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_554_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_554_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_554_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_554_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_554_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_554_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_554_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_555_clock; // @[pe.scala 187:13]
  wire  PE_555_reset; // @[pe.scala 187:13]
  wire  PE_555_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_555_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_555_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_555_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_555_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_555_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_555_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_555_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_555_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_555_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_555_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_556_clock; // @[pe.scala 187:13]
  wire  PE_556_reset; // @[pe.scala 187:13]
  wire  PE_556_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_556_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_556_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_556_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_556_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_556_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_556_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_556_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_556_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_556_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_556_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_557_clock; // @[pe.scala 187:13]
  wire  PE_557_reset; // @[pe.scala 187:13]
  wire  PE_557_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_557_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_557_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_557_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_557_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_557_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_557_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_557_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_557_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_557_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_557_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_558_clock; // @[pe.scala 187:13]
  wire  PE_558_reset; // @[pe.scala 187:13]
  wire  PE_558_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_558_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_558_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_558_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_558_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_558_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_558_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_558_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_558_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_558_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_558_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_559_clock; // @[pe.scala 187:13]
  wire  PE_559_reset; // @[pe.scala 187:13]
  wire  PE_559_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_559_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_559_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_559_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_559_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_559_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_559_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_559_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_559_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_559_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_559_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_560_clock; // @[pe.scala 187:13]
  wire  PE_560_reset; // @[pe.scala 187:13]
  wire  PE_560_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_560_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_560_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_560_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_560_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_560_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_560_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_560_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_560_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_560_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_560_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_561_clock; // @[pe.scala 187:13]
  wire  PE_561_reset; // @[pe.scala 187:13]
  wire  PE_561_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_561_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_561_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_561_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_561_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_561_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_561_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_561_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_561_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_561_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_561_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_562_clock; // @[pe.scala 187:13]
  wire  PE_562_reset; // @[pe.scala 187:13]
  wire  PE_562_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_562_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_562_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_562_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_562_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_562_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_562_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_562_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_562_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_562_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_562_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_563_clock; // @[pe.scala 187:13]
  wire  PE_563_reset; // @[pe.scala 187:13]
  wire  PE_563_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_563_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_563_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_563_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_563_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_563_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_563_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_563_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_563_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_563_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_563_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_564_clock; // @[pe.scala 187:13]
  wire  PE_564_reset; // @[pe.scala 187:13]
  wire  PE_564_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_564_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_564_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_564_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_564_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_564_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_564_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_564_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_564_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_564_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_564_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_565_clock; // @[pe.scala 187:13]
  wire  PE_565_reset; // @[pe.scala 187:13]
  wire  PE_565_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_565_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_565_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_565_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_565_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_565_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_565_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_565_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_565_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_565_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_565_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_566_clock; // @[pe.scala 187:13]
  wire  PE_566_reset; // @[pe.scala 187:13]
  wire  PE_566_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_566_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_566_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_566_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_566_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_566_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_566_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_566_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_566_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_566_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_566_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_567_clock; // @[pe.scala 187:13]
  wire  PE_567_reset; // @[pe.scala 187:13]
  wire  PE_567_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_567_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_567_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_567_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_567_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_567_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_567_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_567_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_567_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_567_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_567_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_568_clock; // @[pe.scala 187:13]
  wire  PE_568_reset; // @[pe.scala 187:13]
  wire  PE_568_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_568_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_568_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_568_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_568_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_568_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_568_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_568_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_568_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_568_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_568_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_569_clock; // @[pe.scala 187:13]
  wire  PE_569_reset; // @[pe.scala 187:13]
  wire  PE_569_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_569_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_569_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_569_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_569_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_569_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_569_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_569_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_569_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_569_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_569_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_570_clock; // @[pe.scala 187:13]
  wire  PE_570_reset; // @[pe.scala 187:13]
  wire  PE_570_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_570_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_570_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_570_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_570_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_570_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_570_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_570_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_570_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_570_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_570_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_571_clock; // @[pe.scala 187:13]
  wire  PE_571_reset; // @[pe.scala 187:13]
  wire  PE_571_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_571_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_571_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_571_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_571_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_571_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_571_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_571_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_571_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_571_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_571_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_572_clock; // @[pe.scala 187:13]
  wire  PE_572_reset; // @[pe.scala 187:13]
  wire  PE_572_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_572_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_572_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_572_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_572_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_572_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_572_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_572_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_572_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_572_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_572_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_573_clock; // @[pe.scala 187:13]
  wire  PE_573_reset; // @[pe.scala 187:13]
  wire  PE_573_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_573_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_573_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_573_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_573_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_573_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_573_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_573_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_573_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_573_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_573_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_574_clock; // @[pe.scala 187:13]
  wire  PE_574_reset; // @[pe.scala 187:13]
  wire  PE_574_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_574_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_574_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_574_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_574_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_574_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_574_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_574_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_574_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_574_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_574_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_575_clock; // @[pe.scala 187:13]
  wire  PE_575_reset; // @[pe.scala 187:13]
  wire  PE_575_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_575_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_575_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_575_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_575_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_575_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_575_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_575_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_575_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_575_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_575_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_576_clock; // @[pe.scala 187:13]
  wire  PE_576_reset; // @[pe.scala 187:13]
  wire  PE_576_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_576_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_576_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_576_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_576_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_576_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_576_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_576_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_576_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_576_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_576_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_577_clock; // @[pe.scala 187:13]
  wire  PE_577_reset; // @[pe.scala 187:13]
  wire  PE_577_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_577_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_577_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_577_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_577_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_577_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_577_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_577_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_577_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_577_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_577_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_578_clock; // @[pe.scala 187:13]
  wire  PE_578_reset; // @[pe.scala 187:13]
  wire  PE_578_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_578_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_578_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_578_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_578_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_578_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_578_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_578_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_578_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_578_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_578_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_579_clock; // @[pe.scala 187:13]
  wire  PE_579_reset; // @[pe.scala 187:13]
  wire  PE_579_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_579_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_579_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_579_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_579_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_579_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_579_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_579_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_579_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_579_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_579_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_580_clock; // @[pe.scala 187:13]
  wire  PE_580_reset; // @[pe.scala 187:13]
  wire  PE_580_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_580_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_580_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_580_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_580_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_580_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_580_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_580_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_580_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_580_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_580_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_581_clock; // @[pe.scala 187:13]
  wire  PE_581_reset; // @[pe.scala 187:13]
  wire  PE_581_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_581_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_581_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_581_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_581_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_581_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_581_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_581_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_581_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_581_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_581_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_582_clock; // @[pe.scala 187:13]
  wire  PE_582_reset; // @[pe.scala 187:13]
  wire  PE_582_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_582_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_582_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_582_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_582_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_582_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_582_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_582_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_582_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_582_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_582_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_583_clock; // @[pe.scala 187:13]
  wire  PE_583_reset; // @[pe.scala 187:13]
  wire  PE_583_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_583_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_583_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_583_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_583_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_583_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_583_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_583_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_583_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_583_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_583_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_584_clock; // @[pe.scala 187:13]
  wire  PE_584_reset; // @[pe.scala 187:13]
  wire  PE_584_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_584_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_584_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_584_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_584_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_584_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_584_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_584_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_584_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_584_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_584_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_585_clock; // @[pe.scala 187:13]
  wire  PE_585_reset; // @[pe.scala 187:13]
  wire  PE_585_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_585_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_585_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_585_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_585_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_585_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_585_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_585_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_585_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_585_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_585_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_586_clock; // @[pe.scala 187:13]
  wire  PE_586_reset; // @[pe.scala 187:13]
  wire  PE_586_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_586_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_586_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_586_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_586_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_586_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_586_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_586_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_586_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_586_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_586_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_587_clock; // @[pe.scala 187:13]
  wire  PE_587_reset; // @[pe.scala 187:13]
  wire  PE_587_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_587_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_587_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_587_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_587_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_587_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_587_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_587_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_587_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_587_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_587_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_588_clock; // @[pe.scala 187:13]
  wire  PE_588_reset; // @[pe.scala 187:13]
  wire  PE_588_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_588_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_588_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_588_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_588_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_588_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_588_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_588_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_588_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_588_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_588_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_589_clock; // @[pe.scala 187:13]
  wire  PE_589_reset; // @[pe.scala 187:13]
  wire  PE_589_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_589_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_589_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_589_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_589_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_589_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_589_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_589_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_589_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_589_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_589_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_590_clock; // @[pe.scala 187:13]
  wire  PE_590_reset; // @[pe.scala 187:13]
  wire  PE_590_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_590_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_590_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_590_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_590_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_590_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_590_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_590_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_590_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_590_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_590_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_591_clock; // @[pe.scala 187:13]
  wire  PE_591_reset; // @[pe.scala 187:13]
  wire  PE_591_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_591_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_591_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_591_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_591_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_591_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_591_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_591_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_591_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_591_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_591_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_592_clock; // @[pe.scala 187:13]
  wire  PE_592_reset; // @[pe.scala 187:13]
  wire  PE_592_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_592_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_592_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_592_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_592_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_592_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_592_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_592_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_592_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_592_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_592_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_593_clock; // @[pe.scala 187:13]
  wire  PE_593_reset; // @[pe.scala 187:13]
  wire  PE_593_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_593_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_593_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_593_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_593_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_593_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_593_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_593_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_593_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_593_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_593_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_594_clock; // @[pe.scala 187:13]
  wire  PE_594_reset; // @[pe.scala 187:13]
  wire  PE_594_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_594_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_594_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_594_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_594_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_594_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_594_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_594_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_594_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_594_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_594_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_595_clock; // @[pe.scala 187:13]
  wire  PE_595_reset; // @[pe.scala 187:13]
  wire  PE_595_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_595_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_595_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_595_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_595_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_595_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_595_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_595_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_595_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_595_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_595_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_596_clock; // @[pe.scala 187:13]
  wire  PE_596_reset; // @[pe.scala 187:13]
  wire  PE_596_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_596_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_596_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_596_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_596_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_596_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_596_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_596_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_596_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_596_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_596_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_597_clock; // @[pe.scala 187:13]
  wire  PE_597_reset; // @[pe.scala 187:13]
  wire  PE_597_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_597_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_597_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_597_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_597_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_597_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_597_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_597_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_597_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_597_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_597_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_598_clock; // @[pe.scala 187:13]
  wire  PE_598_reset; // @[pe.scala 187:13]
  wire  PE_598_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_598_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_598_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_598_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_598_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_598_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_598_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_598_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_598_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_598_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_598_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_599_clock; // @[pe.scala 187:13]
  wire  PE_599_reset; // @[pe.scala 187:13]
  wire  PE_599_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_599_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_599_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_599_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_599_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_599_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_599_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_599_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_599_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_599_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_599_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_600_clock; // @[pe.scala 187:13]
  wire  PE_600_reset; // @[pe.scala 187:13]
  wire  PE_600_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_600_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_600_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_600_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_600_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_600_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_600_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_600_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_600_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_600_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_600_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_601_clock; // @[pe.scala 187:13]
  wire  PE_601_reset; // @[pe.scala 187:13]
  wire  PE_601_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_601_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_601_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_601_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_601_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_601_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_601_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_601_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_601_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_601_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_601_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_602_clock; // @[pe.scala 187:13]
  wire  PE_602_reset; // @[pe.scala 187:13]
  wire  PE_602_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_602_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_602_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_602_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_602_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_602_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_602_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_602_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_602_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_602_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_602_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_603_clock; // @[pe.scala 187:13]
  wire  PE_603_reset; // @[pe.scala 187:13]
  wire  PE_603_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_603_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_603_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_603_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_603_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_603_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_603_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_603_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_603_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_603_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_603_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_604_clock; // @[pe.scala 187:13]
  wire  PE_604_reset; // @[pe.scala 187:13]
  wire  PE_604_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_604_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_604_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_604_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_604_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_604_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_604_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_604_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_604_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_604_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_604_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_605_clock; // @[pe.scala 187:13]
  wire  PE_605_reset; // @[pe.scala 187:13]
  wire  PE_605_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_605_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_605_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_605_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_605_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_605_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_605_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_605_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_605_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_605_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_605_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_606_clock; // @[pe.scala 187:13]
  wire  PE_606_reset; // @[pe.scala 187:13]
  wire  PE_606_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_606_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_606_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_606_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_606_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_606_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_606_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_606_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_606_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_606_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_606_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_607_clock; // @[pe.scala 187:13]
  wire  PE_607_reset; // @[pe.scala 187:13]
  wire  PE_607_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_607_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_607_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_607_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_607_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_607_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_607_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_607_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_607_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_607_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_607_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_608_clock; // @[pe.scala 187:13]
  wire  PE_608_reset; // @[pe.scala 187:13]
  wire  PE_608_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_608_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_608_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_608_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_608_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_608_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_608_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_608_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_608_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_608_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_608_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_609_clock; // @[pe.scala 187:13]
  wire  PE_609_reset; // @[pe.scala 187:13]
  wire  PE_609_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_609_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_609_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_609_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_609_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_609_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_609_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_609_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_609_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_609_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_609_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_610_clock; // @[pe.scala 187:13]
  wire  PE_610_reset; // @[pe.scala 187:13]
  wire  PE_610_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_610_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_610_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_610_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_610_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_610_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_610_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_610_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_610_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_610_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_610_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_611_clock; // @[pe.scala 187:13]
  wire  PE_611_reset; // @[pe.scala 187:13]
  wire  PE_611_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_611_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_611_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_611_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_611_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_611_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_611_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_611_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_611_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_611_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_611_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_612_clock; // @[pe.scala 187:13]
  wire  PE_612_reset; // @[pe.scala 187:13]
  wire  PE_612_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_612_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_612_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_612_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_612_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_612_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_612_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_612_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_612_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_612_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_612_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_613_clock; // @[pe.scala 187:13]
  wire  PE_613_reset; // @[pe.scala 187:13]
  wire  PE_613_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_613_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_613_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_613_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_613_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_613_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_613_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_613_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_613_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_613_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_613_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_614_clock; // @[pe.scala 187:13]
  wire  PE_614_reset; // @[pe.scala 187:13]
  wire  PE_614_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_614_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_614_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_614_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_614_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_614_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_614_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_614_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_614_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_614_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_614_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_615_clock; // @[pe.scala 187:13]
  wire  PE_615_reset; // @[pe.scala 187:13]
  wire  PE_615_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_615_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_615_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_615_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_615_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_615_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_615_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_615_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_615_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_615_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_615_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_616_clock; // @[pe.scala 187:13]
  wire  PE_616_reset; // @[pe.scala 187:13]
  wire  PE_616_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_616_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_616_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_616_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_616_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_616_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_616_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_616_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_616_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_616_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_616_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_617_clock; // @[pe.scala 187:13]
  wire  PE_617_reset; // @[pe.scala 187:13]
  wire  PE_617_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_617_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_617_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_617_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_617_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_617_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_617_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_617_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_617_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_617_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_617_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_618_clock; // @[pe.scala 187:13]
  wire  PE_618_reset; // @[pe.scala 187:13]
  wire  PE_618_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_618_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_618_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_618_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_618_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_618_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_618_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_618_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_618_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_618_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_618_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_619_clock; // @[pe.scala 187:13]
  wire  PE_619_reset; // @[pe.scala 187:13]
  wire  PE_619_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_619_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_619_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_619_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_619_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_619_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_619_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_619_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_619_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_619_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_619_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_620_clock; // @[pe.scala 187:13]
  wire  PE_620_reset; // @[pe.scala 187:13]
  wire  PE_620_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_620_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_620_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_620_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_620_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_620_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_620_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_620_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_620_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_620_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_620_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_621_clock; // @[pe.scala 187:13]
  wire  PE_621_reset; // @[pe.scala 187:13]
  wire  PE_621_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_621_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_621_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_621_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_621_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_621_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_621_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_621_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_621_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_621_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_621_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_622_clock; // @[pe.scala 187:13]
  wire  PE_622_reset; // @[pe.scala 187:13]
  wire  PE_622_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_622_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_622_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_622_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_622_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_622_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_622_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_622_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_622_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_622_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_622_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_623_clock; // @[pe.scala 187:13]
  wire  PE_623_reset; // @[pe.scala 187:13]
  wire  PE_623_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_623_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_623_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_623_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_623_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_623_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_623_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_623_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_623_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_623_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_623_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_624_clock; // @[pe.scala 187:13]
  wire  PE_624_reset; // @[pe.scala 187:13]
  wire  PE_624_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_624_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_624_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_624_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_624_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_624_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_624_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_624_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_624_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_624_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_624_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_625_clock; // @[pe.scala 187:13]
  wire  PE_625_reset; // @[pe.scala 187:13]
  wire  PE_625_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_625_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_625_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_625_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_625_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_625_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_625_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_625_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_625_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_625_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_625_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_626_clock; // @[pe.scala 187:13]
  wire  PE_626_reset; // @[pe.scala 187:13]
  wire  PE_626_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_626_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_626_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_626_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_626_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_626_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_626_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_626_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_626_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_626_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_626_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_627_clock; // @[pe.scala 187:13]
  wire  PE_627_reset; // @[pe.scala 187:13]
  wire  PE_627_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_627_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_627_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_627_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_627_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_627_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_627_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_627_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_627_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_627_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_627_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_628_clock; // @[pe.scala 187:13]
  wire  PE_628_reset; // @[pe.scala 187:13]
  wire  PE_628_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_628_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_628_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_628_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_628_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_628_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_628_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_628_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_628_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_628_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_628_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_629_clock; // @[pe.scala 187:13]
  wire  PE_629_reset; // @[pe.scala 187:13]
  wire  PE_629_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_629_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_629_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_629_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_629_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_629_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_629_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_629_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_629_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_629_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_629_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_630_clock; // @[pe.scala 187:13]
  wire  PE_630_reset; // @[pe.scala 187:13]
  wire  PE_630_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_630_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_630_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_630_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_630_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_630_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_630_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_630_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_630_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_630_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_630_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_631_clock; // @[pe.scala 187:13]
  wire  PE_631_reset; // @[pe.scala 187:13]
  wire  PE_631_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_631_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_631_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_631_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_631_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_631_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_631_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_631_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_631_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_631_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_631_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_632_clock; // @[pe.scala 187:13]
  wire  PE_632_reset; // @[pe.scala 187:13]
  wire  PE_632_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_632_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_632_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_632_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_632_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_632_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_632_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_632_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_632_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_632_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_632_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_633_clock; // @[pe.scala 187:13]
  wire  PE_633_reset; // @[pe.scala 187:13]
  wire  PE_633_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_633_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_633_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_633_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_633_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_633_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_633_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_633_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_633_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_633_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_633_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_634_clock; // @[pe.scala 187:13]
  wire  PE_634_reset; // @[pe.scala 187:13]
  wire  PE_634_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_634_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_634_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_634_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_634_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_634_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_634_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_634_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_634_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_634_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_634_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_635_clock; // @[pe.scala 187:13]
  wire  PE_635_reset; // @[pe.scala 187:13]
  wire  PE_635_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_635_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_635_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_635_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_635_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_635_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_635_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_635_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_635_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_635_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_635_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_636_clock; // @[pe.scala 187:13]
  wire  PE_636_reset; // @[pe.scala 187:13]
  wire  PE_636_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_636_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_636_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_636_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_636_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_636_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_636_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_636_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_636_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_636_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_636_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_637_clock; // @[pe.scala 187:13]
  wire  PE_637_reset; // @[pe.scala 187:13]
  wire  PE_637_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_637_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_637_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_637_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_637_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_637_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_637_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_637_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_637_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_637_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_637_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_638_clock; // @[pe.scala 187:13]
  wire  PE_638_reset; // @[pe.scala 187:13]
  wire  PE_638_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_638_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_638_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_638_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_638_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_638_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_638_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_638_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_638_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_638_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_638_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_639_clock; // @[pe.scala 187:13]
  wire  PE_639_reset; // @[pe.scala 187:13]
  wire  PE_639_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_639_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_639_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_639_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_639_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_639_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_639_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_639_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_639_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_639_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_639_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_640_clock; // @[pe.scala 187:13]
  wire  PE_640_reset; // @[pe.scala 187:13]
  wire  PE_640_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_640_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_640_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_640_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_640_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_640_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_640_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_640_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_640_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_640_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_640_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_641_clock; // @[pe.scala 187:13]
  wire  PE_641_reset; // @[pe.scala 187:13]
  wire  PE_641_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_641_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_641_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_641_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_641_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_641_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_641_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_641_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_641_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_641_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_641_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_642_clock; // @[pe.scala 187:13]
  wire  PE_642_reset; // @[pe.scala 187:13]
  wire  PE_642_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_642_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_642_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_642_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_642_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_642_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_642_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_642_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_642_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_642_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_642_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_643_clock; // @[pe.scala 187:13]
  wire  PE_643_reset; // @[pe.scala 187:13]
  wire  PE_643_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_643_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_643_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_643_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_643_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_643_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_643_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_643_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_643_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_643_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_643_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_644_clock; // @[pe.scala 187:13]
  wire  PE_644_reset; // @[pe.scala 187:13]
  wire  PE_644_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_644_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_644_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_644_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_644_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_644_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_644_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_644_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_644_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_644_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_644_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_645_clock; // @[pe.scala 187:13]
  wire  PE_645_reset; // @[pe.scala 187:13]
  wire  PE_645_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_645_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_645_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_645_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_645_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_645_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_645_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_645_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_645_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_645_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_645_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_646_clock; // @[pe.scala 187:13]
  wire  PE_646_reset; // @[pe.scala 187:13]
  wire  PE_646_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_646_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_646_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_646_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_646_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_646_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_646_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_646_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_646_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_646_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_646_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_647_clock; // @[pe.scala 187:13]
  wire  PE_647_reset; // @[pe.scala 187:13]
  wire  PE_647_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_647_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_647_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_647_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_647_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_647_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_647_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_647_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_647_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_647_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_647_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_648_clock; // @[pe.scala 187:13]
  wire  PE_648_reset; // @[pe.scala 187:13]
  wire  PE_648_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_648_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_648_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_648_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_648_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_648_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_648_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_648_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_648_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_648_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_648_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_649_clock; // @[pe.scala 187:13]
  wire  PE_649_reset; // @[pe.scala 187:13]
  wire  PE_649_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_649_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_649_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_649_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_649_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_649_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_649_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_649_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_649_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_649_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_649_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_650_clock; // @[pe.scala 187:13]
  wire  PE_650_reset; // @[pe.scala 187:13]
  wire  PE_650_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_650_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_650_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_650_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_650_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_650_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_650_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_650_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_650_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_650_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_650_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_651_clock; // @[pe.scala 187:13]
  wire  PE_651_reset; // @[pe.scala 187:13]
  wire  PE_651_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_651_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_651_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_651_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_651_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_651_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_651_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_651_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_651_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_651_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_651_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_652_clock; // @[pe.scala 187:13]
  wire  PE_652_reset; // @[pe.scala 187:13]
  wire  PE_652_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_652_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_652_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_652_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_652_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_652_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_652_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_652_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_652_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_652_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_652_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_653_clock; // @[pe.scala 187:13]
  wire  PE_653_reset; // @[pe.scala 187:13]
  wire  PE_653_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_653_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_653_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_653_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_653_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_653_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_653_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_653_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_653_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_653_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_653_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_654_clock; // @[pe.scala 187:13]
  wire  PE_654_reset; // @[pe.scala 187:13]
  wire  PE_654_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_654_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_654_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_654_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_654_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_654_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_654_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_654_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_654_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_654_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_654_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_655_clock; // @[pe.scala 187:13]
  wire  PE_655_reset; // @[pe.scala 187:13]
  wire  PE_655_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_655_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_655_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_655_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_655_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_655_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_655_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_655_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_655_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_655_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_655_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_656_clock; // @[pe.scala 187:13]
  wire  PE_656_reset; // @[pe.scala 187:13]
  wire  PE_656_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_656_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_656_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_656_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_656_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_656_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_656_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_656_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_656_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_656_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_656_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_657_clock; // @[pe.scala 187:13]
  wire  PE_657_reset; // @[pe.scala 187:13]
  wire  PE_657_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_657_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_657_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_657_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_657_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_657_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_657_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_657_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_657_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_657_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_657_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_658_clock; // @[pe.scala 187:13]
  wire  PE_658_reset; // @[pe.scala 187:13]
  wire  PE_658_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_658_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_658_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_658_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_658_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_658_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_658_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_658_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_658_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_658_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_658_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PE_659_clock; // @[pe.scala 187:13]
  wire  PE_659_reset; // @[pe.scala 187:13]
  wire  PE_659_io_data_2_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_659_io_data_2_out_bits; // @[pe.scala 187:13]
  wire  PE_659_io_data_2_sig_stat2trans; // @[pe.scala 187:13]
  wire  PE_659_io_data_1_in_valid; // @[pe.scala 187:13]
  wire [127:0] PE_659_io_data_1_in_bits; // @[pe.scala 187:13]
  wire  PE_659_io_data_1_out_valid; // @[pe.scala 187:13]
  wire [127:0] PE_659_io_data_1_out_bits; // @[pe.scala 187:13]
  wire  PE_659_io_data_0_in_valid; // @[pe.scala 187:13]
  wire [15:0] PE_659_io_data_0_in_bits; // @[pe.scala 187:13]
  wire  PE_659_io_data_0_out_valid; // @[pe.scala 187:13]
  wire [15:0] PE_659_io_data_0_out_bits; // @[pe.scala 187:13]
  wire  PENetwork_io_to_pes_0_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_io_to_pes_0_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_io_to_pes_1_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_io_to_pes_1_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_io_to_pes_2_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_io_to_pes_2_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_io_to_pes_3_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_io_to_pes_3_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_io_to_pes_4_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_io_to_pes_4_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_io_to_pes_5_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_io_to_pes_5_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_io_to_pes_6_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_io_to_pes_6_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_io_to_pes_7_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_io_to_pes_7_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_io_to_pes_8_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_io_to_pes_8_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_io_to_pes_9_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_io_to_pes_9_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_io_to_pes_10_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_io_to_pes_10_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_io_to_pes_11_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_io_to_pes_11_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_io_to_pes_12_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_io_to_pes_12_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_io_to_pes_13_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_io_to_pes_13_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_io_to_pes_14_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_io_to_pes_14_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_io_to_pes_15_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_io_to_pes_15_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_io_to_pes_16_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_io_to_pes_16_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_io_to_pes_17_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_io_to_pes_17_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_io_to_pes_18_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_io_to_pes_18_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_io_to_pes_19_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_io_to_pes_19_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_io_to_pes_20_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_io_to_pes_20_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_io_to_pes_21_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_io_to_pes_21_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_io_to_pes_21_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_io_to_pes_21_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_io_to_pes_22_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_io_to_pes_22_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_io_to_pes_22_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_io_to_pes_22_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_io_to_pes_23_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_io_to_pes_23_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_io_to_pes_23_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_io_to_pes_23_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_io_to_pes_24_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_io_to_pes_24_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_io_to_pes_24_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_io_to_pes_24_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_io_to_pes_25_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_io_to_pes_25_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_io_to_pes_25_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_io_to_pes_25_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_io_to_pes_26_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_io_to_pes_26_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_io_to_pes_26_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_io_to_pes_26_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_io_to_pes_27_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_io_to_pes_27_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_io_to_pes_27_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_io_to_pes_27_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_io_to_pes_28_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_io_to_pes_28_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_io_to_pes_28_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_io_to_pes_28_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_io_to_pes_29_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_io_to_pes_29_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_io_to_mem_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_1_io_to_pes_0_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_1_io_to_pes_0_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_1_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_1_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_1_io_to_pes_1_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_1_io_to_pes_1_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_1_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_1_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_1_io_to_pes_2_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_1_io_to_pes_2_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_1_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_1_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_1_io_to_pes_3_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_1_io_to_pes_3_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_1_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_1_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_1_io_to_pes_4_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_1_io_to_pes_4_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_1_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_1_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_1_io_to_pes_5_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_1_io_to_pes_5_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_1_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_1_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_1_io_to_pes_6_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_1_io_to_pes_6_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_1_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_1_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_1_io_to_pes_7_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_1_io_to_pes_7_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_1_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_1_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_1_io_to_pes_8_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_1_io_to_pes_8_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_1_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_1_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_1_io_to_pes_9_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_1_io_to_pes_9_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_1_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_1_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_1_io_to_pes_10_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_1_io_to_pes_10_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_1_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_1_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_1_io_to_pes_11_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_1_io_to_pes_11_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_1_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_1_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_1_io_to_pes_12_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_1_io_to_pes_12_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_1_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_1_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_1_io_to_pes_13_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_1_io_to_pes_13_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_1_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_1_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_1_io_to_pes_14_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_1_io_to_pes_14_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_1_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_1_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_1_io_to_pes_15_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_1_io_to_pes_15_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_1_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_1_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_1_io_to_pes_16_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_1_io_to_pes_16_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_1_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_1_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_1_io_to_pes_17_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_1_io_to_pes_17_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_1_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_1_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_1_io_to_pes_18_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_1_io_to_pes_18_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_1_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_1_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_1_io_to_pes_19_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_1_io_to_pes_19_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_1_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_1_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_1_io_to_pes_20_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_1_io_to_pes_20_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_1_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_1_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_1_io_to_pes_21_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_1_io_to_pes_21_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_1_io_to_pes_21_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_1_io_to_pes_21_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_1_io_to_pes_22_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_1_io_to_pes_22_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_1_io_to_pes_22_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_1_io_to_pes_22_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_1_io_to_pes_23_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_1_io_to_pes_23_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_1_io_to_pes_23_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_1_io_to_pes_23_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_1_io_to_pes_24_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_1_io_to_pes_24_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_1_io_to_pes_24_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_1_io_to_pes_24_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_1_io_to_pes_25_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_1_io_to_pes_25_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_1_io_to_pes_25_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_1_io_to_pes_25_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_1_io_to_pes_26_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_1_io_to_pes_26_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_1_io_to_pes_26_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_1_io_to_pes_26_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_1_io_to_pes_27_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_1_io_to_pes_27_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_1_io_to_pes_27_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_1_io_to_pes_27_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_1_io_to_pes_28_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_1_io_to_pes_28_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_1_io_to_pes_28_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_1_io_to_pes_28_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_1_io_to_pes_29_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_1_io_to_pes_29_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_1_io_to_mem_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_1_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_2_io_to_pes_0_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_2_io_to_pes_0_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_2_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_2_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_2_io_to_pes_1_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_2_io_to_pes_1_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_2_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_2_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_2_io_to_pes_2_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_2_io_to_pes_2_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_2_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_2_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_2_io_to_pes_3_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_2_io_to_pes_3_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_2_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_2_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_2_io_to_pes_4_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_2_io_to_pes_4_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_2_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_2_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_2_io_to_pes_5_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_2_io_to_pes_5_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_2_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_2_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_2_io_to_pes_6_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_2_io_to_pes_6_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_2_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_2_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_2_io_to_pes_7_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_2_io_to_pes_7_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_2_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_2_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_2_io_to_pes_8_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_2_io_to_pes_8_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_2_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_2_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_2_io_to_pes_9_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_2_io_to_pes_9_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_2_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_2_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_2_io_to_pes_10_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_2_io_to_pes_10_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_2_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_2_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_2_io_to_pes_11_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_2_io_to_pes_11_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_2_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_2_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_2_io_to_pes_12_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_2_io_to_pes_12_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_2_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_2_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_2_io_to_pes_13_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_2_io_to_pes_13_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_2_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_2_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_2_io_to_pes_14_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_2_io_to_pes_14_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_2_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_2_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_2_io_to_pes_15_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_2_io_to_pes_15_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_2_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_2_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_2_io_to_pes_16_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_2_io_to_pes_16_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_2_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_2_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_2_io_to_pes_17_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_2_io_to_pes_17_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_2_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_2_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_2_io_to_pes_18_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_2_io_to_pes_18_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_2_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_2_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_2_io_to_pes_19_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_2_io_to_pes_19_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_2_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_2_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_2_io_to_pes_20_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_2_io_to_pes_20_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_2_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_2_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_2_io_to_pes_21_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_2_io_to_pes_21_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_2_io_to_pes_21_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_2_io_to_pes_21_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_2_io_to_pes_22_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_2_io_to_pes_22_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_2_io_to_pes_22_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_2_io_to_pes_22_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_2_io_to_pes_23_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_2_io_to_pes_23_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_2_io_to_pes_23_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_2_io_to_pes_23_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_2_io_to_pes_24_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_2_io_to_pes_24_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_2_io_to_pes_24_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_2_io_to_pes_24_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_2_io_to_pes_25_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_2_io_to_pes_25_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_2_io_to_pes_25_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_2_io_to_pes_25_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_2_io_to_pes_26_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_2_io_to_pes_26_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_2_io_to_pes_26_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_2_io_to_pes_26_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_2_io_to_pes_27_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_2_io_to_pes_27_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_2_io_to_pes_27_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_2_io_to_pes_27_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_2_io_to_pes_28_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_2_io_to_pes_28_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_2_io_to_pes_28_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_2_io_to_pes_28_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_2_io_to_pes_29_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_2_io_to_pes_29_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_2_io_to_mem_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_2_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_3_io_to_pes_0_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_3_io_to_pes_0_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_3_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_3_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_3_io_to_pes_1_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_3_io_to_pes_1_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_3_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_3_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_3_io_to_pes_2_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_3_io_to_pes_2_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_3_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_3_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_3_io_to_pes_3_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_3_io_to_pes_3_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_3_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_3_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_3_io_to_pes_4_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_3_io_to_pes_4_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_3_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_3_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_3_io_to_pes_5_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_3_io_to_pes_5_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_3_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_3_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_3_io_to_pes_6_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_3_io_to_pes_6_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_3_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_3_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_3_io_to_pes_7_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_3_io_to_pes_7_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_3_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_3_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_3_io_to_pes_8_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_3_io_to_pes_8_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_3_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_3_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_3_io_to_pes_9_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_3_io_to_pes_9_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_3_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_3_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_3_io_to_pes_10_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_3_io_to_pes_10_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_3_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_3_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_3_io_to_pes_11_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_3_io_to_pes_11_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_3_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_3_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_3_io_to_pes_12_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_3_io_to_pes_12_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_3_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_3_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_3_io_to_pes_13_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_3_io_to_pes_13_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_3_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_3_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_3_io_to_pes_14_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_3_io_to_pes_14_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_3_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_3_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_3_io_to_pes_15_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_3_io_to_pes_15_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_3_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_3_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_3_io_to_pes_16_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_3_io_to_pes_16_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_3_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_3_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_3_io_to_pes_17_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_3_io_to_pes_17_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_3_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_3_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_3_io_to_pes_18_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_3_io_to_pes_18_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_3_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_3_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_3_io_to_pes_19_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_3_io_to_pes_19_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_3_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_3_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_3_io_to_pes_20_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_3_io_to_pes_20_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_3_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_3_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_3_io_to_pes_21_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_3_io_to_pes_21_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_3_io_to_pes_21_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_3_io_to_pes_21_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_3_io_to_pes_22_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_3_io_to_pes_22_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_3_io_to_pes_22_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_3_io_to_pes_22_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_3_io_to_pes_23_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_3_io_to_pes_23_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_3_io_to_pes_23_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_3_io_to_pes_23_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_3_io_to_pes_24_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_3_io_to_pes_24_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_3_io_to_pes_24_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_3_io_to_pes_24_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_3_io_to_pes_25_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_3_io_to_pes_25_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_3_io_to_pes_25_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_3_io_to_pes_25_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_3_io_to_pes_26_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_3_io_to_pes_26_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_3_io_to_pes_26_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_3_io_to_pes_26_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_3_io_to_pes_27_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_3_io_to_pes_27_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_3_io_to_pes_27_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_3_io_to_pes_27_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_3_io_to_pes_28_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_3_io_to_pes_28_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_3_io_to_pes_28_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_3_io_to_pes_28_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_3_io_to_pes_29_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_3_io_to_pes_29_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_3_io_to_mem_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_3_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_4_io_to_pes_0_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_4_io_to_pes_0_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_4_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_4_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_4_io_to_pes_1_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_4_io_to_pes_1_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_4_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_4_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_4_io_to_pes_2_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_4_io_to_pes_2_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_4_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_4_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_4_io_to_pes_3_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_4_io_to_pes_3_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_4_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_4_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_4_io_to_pes_4_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_4_io_to_pes_4_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_4_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_4_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_4_io_to_pes_5_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_4_io_to_pes_5_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_4_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_4_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_4_io_to_pes_6_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_4_io_to_pes_6_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_4_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_4_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_4_io_to_pes_7_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_4_io_to_pes_7_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_4_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_4_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_4_io_to_pes_8_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_4_io_to_pes_8_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_4_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_4_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_4_io_to_pes_9_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_4_io_to_pes_9_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_4_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_4_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_4_io_to_pes_10_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_4_io_to_pes_10_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_4_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_4_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_4_io_to_pes_11_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_4_io_to_pes_11_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_4_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_4_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_4_io_to_pes_12_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_4_io_to_pes_12_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_4_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_4_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_4_io_to_pes_13_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_4_io_to_pes_13_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_4_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_4_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_4_io_to_pes_14_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_4_io_to_pes_14_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_4_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_4_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_4_io_to_pes_15_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_4_io_to_pes_15_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_4_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_4_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_4_io_to_pes_16_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_4_io_to_pes_16_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_4_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_4_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_4_io_to_pes_17_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_4_io_to_pes_17_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_4_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_4_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_4_io_to_pes_18_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_4_io_to_pes_18_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_4_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_4_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_4_io_to_pes_19_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_4_io_to_pes_19_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_4_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_4_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_4_io_to_pes_20_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_4_io_to_pes_20_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_4_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_4_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_4_io_to_pes_21_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_4_io_to_pes_21_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_4_io_to_pes_21_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_4_io_to_pes_21_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_4_io_to_pes_22_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_4_io_to_pes_22_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_4_io_to_pes_22_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_4_io_to_pes_22_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_4_io_to_pes_23_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_4_io_to_pes_23_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_4_io_to_pes_23_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_4_io_to_pes_23_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_4_io_to_pes_24_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_4_io_to_pes_24_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_4_io_to_pes_24_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_4_io_to_pes_24_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_4_io_to_pes_25_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_4_io_to_pes_25_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_4_io_to_pes_25_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_4_io_to_pes_25_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_4_io_to_pes_26_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_4_io_to_pes_26_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_4_io_to_pes_26_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_4_io_to_pes_26_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_4_io_to_pes_27_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_4_io_to_pes_27_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_4_io_to_pes_27_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_4_io_to_pes_27_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_4_io_to_pes_28_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_4_io_to_pes_28_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_4_io_to_pes_28_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_4_io_to_pes_28_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_4_io_to_pes_29_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_4_io_to_pes_29_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_4_io_to_mem_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_4_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_5_io_to_pes_0_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_5_io_to_pes_0_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_5_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_5_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_5_io_to_pes_1_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_5_io_to_pes_1_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_5_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_5_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_5_io_to_pes_2_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_5_io_to_pes_2_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_5_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_5_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_5_io_to_pes_3_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_5_io_to_pes_3_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_5_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_5_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_5_io_to_pes_4_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_5_io_to_pes_4_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_5_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_5_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_5_io_to_pes_5_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_5_io_to_pes_5_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_5_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_5_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_5_io_to_pes_6_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_5_io_to_pes_6_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_5_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_5_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_5_io_to_pes_7_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_5_io_to_pes_7_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_5_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_5_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_5_io_to_pes_8_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_5_io_to_pes_8_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_5_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_5_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_5_io_to_pes_9_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_5_io_to_pes_9_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_5_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_5_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_5_io_to_pes_10_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_5_io_to_pes_10_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_5_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_5_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_5_io_to_pes_11_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_5_io_to_pes_11_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_5_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_5_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_5_io_to_pes_12_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_5_io_to_pes_12_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_5_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_5_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_5_io_to_pes_13_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_5_io_to_pes_13_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_5_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_5_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_5_io_to_pes_14_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_5_io_to_pes_14_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_5_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_5_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_5_io_to_pes_15_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_5_io_to_pes_15_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_5_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_5_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_5_io_to_pes_16_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_5_io_to_pes_16_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_5_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_5_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_5_io_to_pes_17_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_5_io_to_pes_17_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_5_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_5_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_5_io_to_pes_18_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_5_io_to_pes_18_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_5_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_5_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_5_io_to_pes_19_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_5_io_to_pes_19_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_5_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_5_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_5_io_to_pes_20_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_5_io_to_pes_20_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_5_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_5_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_5_io_to_pes_21_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_5_io_to_pes_21_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_5_io_to_pes_21_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_5_io_to_pes_21_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_5_io_to_pes_22_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_5_io_to_pes_22_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_5_io_to_pes_22_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_5_io_to_pes_22_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_5_io_to_pes_23_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_5_io_to_pes_23_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_5_io_to_pes_23_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_5_io_to_pes_23_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_5_io_to_pes_24_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_5_io_to_pes_24_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_5_io_to_pes_24_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_5_io_to_pes_24_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_5_io_to_pes_25_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_5_io_to_pes_25_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_5_io_to_pes_25_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_5_io_to_pes_25_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_5_io_to_pes_26_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_5_io_to_pes_26_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_5_io_to_pes_26_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_5_io_to_pes_26_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_5_io_to_pes_27_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_5_io_to_pes_27_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_5_io_to_pes_27_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_5_io_to_pes_27_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_5_io_to_pes_28_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_5_io_to_pes_28_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_5_io_to_pes_28_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_5_io_to_pes_28_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_5_io_to_pes_29_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_5_io_to_pes_29_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_5_io_to_mem_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_5_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_6_io_to_pes_0_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_6_io_to_pes_0_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_6_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_6_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_6_io_to_pes_1_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_6_io_to_pes_1_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_6_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_6_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_6_io_to_pes_2_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_6_io_to_pes_2_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_6_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_6_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_6_io_to_pes_3_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_6_io_to_pes_3_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_6_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_6_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_6_io_to_pes_4_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_6_io_to_pes_4_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_6_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_6_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_6_io_to_pes_5_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_6_io_to_pes_5_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_6_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_6_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_6_io_to_pes_6_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_6_io_to_pes_6_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_6_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_6_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_6_io_to_pes_7_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_6_io_to_pes_7_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_6_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_6_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_6_io_to_pes_8_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_6_io_to_pes_8_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_6_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_6_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_6_io_to_pes_9_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_6_io_to_pes_9_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_6_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_6_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_6_io_to_pes_10_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_6_io_to_pes_10_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_6_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_6_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_6_io_to_pes_11_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_6_io_to_pes_11_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_6_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_6_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_6_io_to_pes_12_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_6_io_to_pes_12_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_6_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_6_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_6_io_to_pes_13_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_6_io_to_pes_13_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_6_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_6_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_6_io_to_pes_14_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_6_io_to_pes_14_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_6_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_6_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_6_io_to_pes_15_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_6_io_to_pes_15_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_6_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_6_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_6_io_to_pes_16_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_6_io_to_pes_16_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_6_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_6_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_6_io_to_pes_17_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_6_io_to_pes_17_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_6_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_6_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_6_io_to_pes_18_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_6_io_to_pes_18_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_6_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_6_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_6_io_to_pes_19_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_6_io_to_pes_19_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_6_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_6_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_6_io_to_pes_20_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_6_io_to_pes_20_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_6_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_6_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_6_io_to_pes_21_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_6_io_to_pes_21_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_6_io_to_pes_21_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_6_io_to_pes_21_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_6_io_to_pes_22_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_6_io_to_pes_22_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_6_io_to_pes_22_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_6_io_to_pes_22_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_6_io_to_pes_23_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_6_io_to_pes_23_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_6_io_to_pes_23_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_6_io_to_pes_23_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_6_io_to_pes_24_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_6_io_to_pes_24_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_6_io_to_pes_24_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_6_io_to_pes_24_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_6_io_to_pes_25_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_6_io_to_pes_25_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_6_io_to_pes_25_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_6_io_to_pes_25_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_6_io_to_pes_26_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_6_io_to_pes_26_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_6_io_to_pes_26_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_6_io_to_pes_26_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_6_io_to_pes_27_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_6_io_to_pes_27_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_6_io_to_pes_27_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_6_io_to_pes_27_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_6_io_to_pes_28_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_6_io_to_pes_28_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_6_io_to_pes_28_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_6_io_to_pes_28_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_6_io_to_pes_29_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_6_io_to_pes_29_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_6_io_to_mem_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_6_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_7_io_to_pes_0_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_7_io_to_pes_0_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_7_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_7_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_7_io_to_pes_1_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_7_io_to_pes_1_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_7_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_7_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_7_io_to_pes_2_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_7_io_to_pes_2_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_7_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_7_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_7_io_to_pes_3_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_7_io_to_pes_3_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_7_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_7_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_7_io_to_pes_4_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_7_io_to_pes_4_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_7_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_7_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_7_io_to_pes_5_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_7_io_to_pes_5_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_7_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_7_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_7_io_to_pes_6_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_7_io_to_pes_6_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_7_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_7_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_7_io_to_pes_7_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_7_io_to_pes_7_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_7_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_7_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_7_io_to_pes_8_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_7_io_to_pes_8_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_7_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_7_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_7_io_to_pes_9_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_7_io_to_pes_9_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_7_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_7_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_7_io_to_pes_10_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_7_io_to_pes_10_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_7_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_7_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_7_io_to_pes_11_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_7_io_to_pes_11_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_7_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_7_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_7_io_to_pes_12_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_7_io_to_pes_12_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_7_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_7_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_7_io_to_pes_13_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_7_io_to_pes_13_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_7_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_7_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_7_io_to_pes_14_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_7_io_to_pes_14_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_7_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_7_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_7_io_to_pes_15_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_7_io_to_pes_15_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_7_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_7_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_7_io_to_pes_16_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_7_io_to_pes_16_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_7_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_7_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_7_io_to_pes_17_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_7_io_to_pes_17_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_7_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_7_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_7_io_to_pes_18_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_7_io_to_pes_18_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_7_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_7_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_7_io_to_pes_19_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_7_io_to_pes_19_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_7_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_7_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_7_io_to_pes_20_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_7_io_to_pes_20_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_7_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_7_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_7_io_to_pes_21_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_7_io_to_pes_21_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_7_io_to_pes_21_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_7_io_to_pes_21_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_7_io_to_pes_22_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_7_io_to_pes_22_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_7_io_to_pes_22_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_7_io_to_pes_22_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_7_io_to_pes_23_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_7_io_to_pes_23_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_7_io_to_pes_23_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_7_io_to_pes_23_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_7_io_to_pes_24_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_7_io_to_pes_24_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_7_io_to_pes_24_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_7_io_to_pes_24_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_7_io_to_pes_25_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_7_io_to_pes_25_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_7_io_to_pes_25_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_7_io_to_pes_25_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_7_io_to_pes_26_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_7_io_to_pes_26_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_7_io_to_pes_26_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_7_io_to_pes_26_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_7_io_to_pes_27_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_7_io_to_pes_27_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_7_io_to_pes_27_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_7_io_to_pes_27_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_7_io_to_pes_28_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_7_io_to_pes_28_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_7_io_to_pes_28_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_7_io_to_pes_28_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_7_io_to_pes_29_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_7_io_to_pes_29_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_7_io_to_mem_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_7_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_8_io_to_pes_0_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_8_io_to_pes_0_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_8_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_8_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_8_io_to_pes_1_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_8_io_to_pes_1_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_8_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_8_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_8_io_to_pes_2_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_8_io_to_pes_2_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_8_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_8_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_8_io_to_pes_3_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_8_io_to_pes_3_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_8_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_8_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_8_io_to_pes_4_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_8_io_to_pes_4_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_8_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_8_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_8_io_to_pes_5_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_8_io_to_pes_5_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_8_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_8_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_8_io_to_pes_6_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_8_io_to_pes_6_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_8_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_8_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_8_io_to_pes_7_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_8_io_to_pes_7_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_8_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_8_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_8_io_to_pes_8_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_8_io_to_pes_8_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_8_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_8_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_8_io_to_pes_9_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_8_io_to_pes_9_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_8_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_8_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_8_io_to_pes_10_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_8_io_to_pes_10_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_8_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_8_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_8_io_to_pes_11_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_8_io_to_pes_11_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_8_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_8_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_8_io_to_pes_12_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_8_io_to_pes_12_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_8_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_8_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_8_io_to_pes_13_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_8_io_to_pes_13_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_8_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_8_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_8_io_to_pes_14_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_8_io_to_pes_14_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_8_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_8_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_8_io_to_pes_15_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_8_io_to_pes_15_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_8_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_8_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_8_io_to_pes_16_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_8_io_to_pes_16_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_8_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_8_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_8_io_to_pes_17_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_8_io_to_pes_17_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_8_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_8_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_8_io_to_pes_18_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_8_io_to_pes_18_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_8_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_8_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_8_io_to_pes_19_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_8_io_to_pes_19_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_8_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_8_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_8_io_to_pes_20_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_8_io_to_pes_20_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_8_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_8_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_8_io_to_pes_21_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_8_io_to_pes_21_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_8_io_to_pes_21_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_8_io_to_pes_21_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_8_io_to_pes_22_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_8_io_to_pes_22_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_8_io_to_pes_22_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_8_io_to_pes_22_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_8_io_to_pes_23_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_8_io_to_pes_23_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_8_io_to_pes_23_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_8_io_to_pes_23_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_8_io_to_pes_24_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_8_io_to_pes_24_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_8_io_to_pes_24_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_8_io_to_pes_24_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_8_io_to_pes_25_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_8_io_to_pes_25_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_8_io_to_pes_25_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_8_io_to_pes_25_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_8_io_to_pes_26_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_8_io_to_pes_26_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_8_io_to_pes_26_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_8_io_to_pes_26_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_8_io_to_pes_27_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_8_io_to_pes_27_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_8_io_to_pes_27_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_8_io_to_pes_27_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_8_io_to_pes_28_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_8_io_to_pes_28_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_8_io_to_pes_28_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_8_io_to_pes_28_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_8_io_to_pes_29_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_8_io_to_pes_29_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_8_io_to_mem_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_8_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_9_io_to_pes_0_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_9_io_to_pes_0_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_9_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_9_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_9_io_to_pes_1_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_9_io_to_pes_1_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_9_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_9_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_9_io_to_pes_2_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_9_io_to_pes_2_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_9_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_9_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_9_io_to_pes_3_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_9_io_to_pes_3_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_9_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_9_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_9_io_to_pes_4_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_9_io_to_pes_4_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_9_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_9_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_9_io_to_pes_5_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_9_io_to_pes_5_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_9_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_9_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_9_io_to_pes_6_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_9_io_to_pes_6_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_9_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_9_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_9_io_to_pes_7_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_9_io_to_pes_7_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_9_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_9_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_9_io_to_pes_8_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_9_io_to_pes_8_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_9_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_9_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_9_io_to_pes_9_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_9_io_to_pes_9_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_9_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_9_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_9_io_to_pes_10_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_9_io_to_pes_10_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_9_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_9_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_9_io_to_pes_11_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_9_io_to_pes_11_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_9_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_9_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_9_io_to_pes_12_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_9_io_to_pes_12_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_9_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_9_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_9_io_to_pes_13_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_9_io_to_pes_13_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_9_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_9_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_9_io_to_pes_14_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_9_io_to_pes_14_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_9_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_9_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_9_io_to_pes_15_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_9_io_to_pes_15_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_9_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_9_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_9_io_to_pes_16_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_9_io_to_pes_16_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_9_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_9_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_9_io_to_pes_17_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_9_io_to_pes_17_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_9_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_9_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_9_io_to_pes_18_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_9_io_to_pes_18_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_9_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_9_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_9_io_to_pes_19_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_9_io_to_pes_19_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_9_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_9_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_9_io_to_pes_20_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_9_io_to_pes_20_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_9_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_9_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_9_io_to_pes_21_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_9_io_to_pes_21_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_9_io_to_pes_21_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_9_io_to_pes_21_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_9_io_to_pes_22_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_9_io_to_pes_22_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_9_io_to_pes_22_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_9_io_to_pes_22_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_9_io_to_pes_23_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_9_io_to_pes_23_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_9_io_to_pes_23_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_9_io_to_pes_23_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_9_io_to_pes_24_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_9_io_to_pes_24_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_9_io_to_pes_24_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_9_io_to_pes_24_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_9_io_to_pes_25_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_9_io_to_pes_25_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_9_io_to_pes_25_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_9_io_to_pes_25_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_9_io_to_pes_26_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_9_io_to_pes_26_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_9_io_to_pes_26_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_9_io_to_pes_26_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_9_io_to_pes_27_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_9_io_to_pes_27_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_9_io_to_pes_27_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_9_io_to_pes_27_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_9_io_to_pes_28_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_9_io_to_pes_28_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_9_io_to_pes_28_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_9_io_to_pes_28_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_9_io_to_pes_29_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_9_io_to_pes_29_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_9_io_to_mem_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_9_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_10_io_to_pes_0_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_10_io_to_pes_0_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_10_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_10_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_10_io_to_pes_1_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_10_io_to_pes_1_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_10_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_10_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_10_io_to_pes_2_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_10_io_to_pes_2_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_10_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_10_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_10_io_to_pes_3_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_10_io_to_pes_3_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_10_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_10_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_10_io_to_pes_4_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_10_io_to_pes_4_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_10_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_10_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_10_io_to_pes_5_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_10_io_to_pes_5_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_10_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_10_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_10_io_to_pes_6_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_10_io_to_pes_6_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_10_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_10_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_10_io_to_pes_7_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_10_io_to_pes_7_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_10_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_10_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_10_io_to_pes_8_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_10_io_to_pes_8_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_10_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_10_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_10_io_to_pes_9_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_10_io_to_pes_9_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_10_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_10_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_10_io_to_pes_10_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_10_io_to_pes_10_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_10_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_10_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_10_io_to_pes_11_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_10_io_to_pes_11_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_10_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_10_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_10_io_to_pes_12_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_10_io_to_pes_12_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_10_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_10_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_10_io_to_pes_13_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_10_io_to_pes_13_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_10_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_10_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_10_io_to_pes_14_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_10_io_to_pes_14_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_10_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_10_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_10_io_to_pes_15_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_10_io_to_pes_15_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_10_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_10_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_10_io_to_pes_16_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_10_io_to_pes_16_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_10_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_10_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_10_io_to_pes_17_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_10_io_to_pes_17_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_10_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_10_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_10_io_to_pes_18_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_10_io_to_pes_18_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_10_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_10_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_10_io_to_pes_19_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_10_io_to_pes_19_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_10_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_10_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_10_io_to_pes_20_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_10_io_to_pes_20_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_10_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_10_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_10_io_to_pes_21_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_10_io_to_pes_21_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_10_io_to_pes_21_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_10_io_to_pes_21_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_10_io_to_pes_22_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_10_io_to_pes_22_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_10_io_to_pes_22_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_10_io_to_pes_22_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_10_io_to_pes_23_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_10_io_to_pes_23_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_10_io_to_pes_23_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_10_io_to_pes_23_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_10_io_to_pes_24_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_10_io_to_pes_24_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_10_io_to_pes_24_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_10_io_to_pes_24_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_10_io_to_pes_25_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_10_io_to_pes_25_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_10_io_to_pes_25_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_10_io_to_pes_25_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_10_io_to_pes_26_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_10_io_to_pes_26_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_10_io_to_pes_26_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_10_io_to_pes_26_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_10_io_to_pes_27_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_10_io_to_pes_27_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_10_io_to_pes_27_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_10_io_to_pes_27_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_10_io_to_pes_28_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_10_io_to_pes_28_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_10_io_to_pes_28_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_10_io_to_pes_28_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_10_io_to_pes_29_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_10_io_to_pes_29_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_10_io_to_mem_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_10_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_11_io_to_pes_0_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_11_io_to_pes_0_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_11_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_11_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_11_io_to_pes_1_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_11_io_to_pes_1_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_11_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_11_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_11_io_to_pes_2_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_11_io_to_pes_2_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_11_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_11_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_11_io_to_pes_3_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_11_io_to_pes_3_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_11_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_11_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_11_io_to_pes_4_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_11_io_to_pes_4_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_11_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_11_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_11_io_to_pes_5_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_11_io_to_pes_5_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_11_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_11_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_11_io_to_pes_6_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_11_io_to_pes_6_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_11_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_11_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_11_io_to_pes_7_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_11_io_to_pes_7_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_11_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_11_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_11_io_to_pes_8_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_11_io_to_pes_8_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_11_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_11_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_11_io_to_pes_9_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_11_io_to_pes_9_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_11_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_11_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_11_io_to_pes_10_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_11_io_to_pes_10_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_11_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_11_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_11_io_to_pes_11_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_11_io_to_pes_11_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_11_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_11_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_11_io_to_pes_12_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_11_io_to_pes_12_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_11_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_11_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_11_io_to_pes_13_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_11_io_to_pes_13_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_11_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_11_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_11_io_to_pes_14_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_11_io_to_pes_14_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_11_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_11_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_11_io_to_pes_15_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_11_io_to_pes_15_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_11_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_11_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_11_io_to_pes_16_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_11_io_to_pes_16_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_11_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_11_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_11_io_to_pes_17_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_11_io_to_pes_17_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_11_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_11_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_11_io_to_pes_18_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_11_io_to_pes_18_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_11_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_11_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_11_io_to_pes_19_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_11_io_to_pes_19_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_11_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_11_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_11_io_to_pes_20_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_11_io_to_pes_20_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_11_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_11_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_11_io_to_pes_21_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_11_io_to_pes_21_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_11_io_to_pes_21_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_11_io_to_pes_21_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_11_io_to_pes_22_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_11_io_to_pes_22_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_11_io_to_pes_22_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_11_io_to_pes_22_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_11_io_to_pes_23_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_11_io_to_pes_23_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_11_io_to_pes_23_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_11_io_to_pes_23_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_11_io_to_pes_24_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_11_io_to_pes_24_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_11_io_to_pes_24_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_11_io_to_pes_24_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_11_io_to_pes_25_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_11_io_to_pes_25_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_11_io_to_pes_25_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_11_io_to_pes_25_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_11_io_to_pes_26_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_11_io_to_pes_26_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_11_io_to_pes_26_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_11_io_to_pes_26_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_11_io_to_pes_27_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_11_io_to_pes_27_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_11_io_to_pes_27_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_11_io_to_pes_27_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_11_io_to_pes_28_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_11_io_to_pes_28_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_11_io_to_pes_28_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_11_io_to_pes_28_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_11_io_to_pes_29_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_11_io_to_pes_29_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_11_io_to_mem_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_11_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_12_io_to_pes_0_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_12_io_to_pes_0_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_12_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_12_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_12_io_to_pes_1_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_12_io_to_pes_1_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_12_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_12_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_12_io_to_pes_2_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_12_io_to_pes_2_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_12_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_12_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_12_io_to_pes_3_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_12_io_to_pes_3_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_12_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_12_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_12_io_to_pes_4_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_12_io_to_pes_4_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_12_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_12_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_12_io_to_pes_5_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_12_io_to_pes_5_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_12_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_12_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_12_io_to_pes_6_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_12_io_to_pes_6_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_12_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_12_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_12_io_to_pes_7_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_12_io_to_pes_7_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_12_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_12_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_12_io_to_pes_8_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_12_io_to_pes_8_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_12_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_12_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_12_io_to_pes_9_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_12_io_to_pes_9_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_12_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_12_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_12_io_to_pes_10_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_12_io_to_pes_10_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_12_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_12_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_12_io_to_pes_11_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_12_io_to_pes_11_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_12_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_12_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_12_io_to_pes_12_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_12_io_to_pes_12_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_12_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_12_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_12_io_to_pes_13_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_12_io_to_pes_13_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_12_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_12_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_12_io_to_pes_14_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_12_io_to_pes_14_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_12_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_12_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_12_io_to_pes_15_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_12_io_to_pes_15_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_12_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_12_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_12_io_to_pes_16_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_12_io_to_pes_16_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_12_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_12_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_12_io_to_pes_17_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_12_io_to_pes_17_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_12_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_12_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_12_io_to_pes_18_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_12_io_to_pes_18_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_12_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_12_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_12_io_to_pes_19_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_12_io_to_pes_19_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_12_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_12_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_12_io_to_pes_20_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_12_io_to_pes_20_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_12_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_12_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_12_io_to_pes_21_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_12_io_to_pes_21_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_12_io_to_pes_21_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_12_io_to_pes_21_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_12_io_to_pes_22_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_12_io_to_pes_22_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_12_io_to_pes_22_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_12_io_to_pes_22_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_12_io_to_pes_23_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_12_io_to_pes_23_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_12_io_to_pes_23_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_12_io_to_pes_23_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_12_io_to_pes_24_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_12_io_to_pes_24_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_12_io_to_pes_24_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_12_io_to_pes_24_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_12_io_to_pes_25_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_12_io_to_pes_25_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_12_io_to_pes_25_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_12_io_to_pes_25_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_12_io_to_pes_26_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_12_io_to_pes_26_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_12_io_to_pes_26_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_12_io_to_pes_26_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_12_io_to_pes_27_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_12_io_to_pes_27_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_12_io_to_pes_27_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_12_io_to_pes_27_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_12_io_to_pes_28_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_12_io_to_pes_28_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_12_io_to_pes_28_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_12_io_to_pes_28_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_12_io_to_pes_29_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_12_io_to_pes_29_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_12_io_to_mem_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_12_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_13_io_to_pes_0_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_13_io_to_pes_0_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_13_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_13_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_13_io_to_pes_1_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_13_io_to_pes_1_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_13_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_13_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_13_io_to_pes_2_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_13_io_to_pes_2_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_13_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_13_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_13_io_to_pes_3_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_13_io_to_pes_3_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_13_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_13_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_13_io_to_pes_4_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_13_io_to_pes_4_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_13_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_13_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_13_io_to_pes_5_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_13_io_to_pes_5_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_13_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_13_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_13_io_to_pes_6_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_13_io_to_pes_6_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_13_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_13_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_13_io_to_pes_7_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_13_io_to_pes_7_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_13_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_13_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_13_io_to_pes_8_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_13_io_to_pes_8_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_13_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_13_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_13_io_to_pes_9_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_13_io_to_pes_9_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_13_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_13_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_13_io_to_pes_10_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_13_io_to_pes_10_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_13_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_13_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_13_io_to_pes_11_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_13_io_to_pes_11_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_13_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_13_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_13_io_to_pes_12_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_13_io_to_pes_12_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_13_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_13_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_13_io_to_pes_13_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_13_io_to_pes_13_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_13_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_13_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_13_io_to_pes_14_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_13_io_to_pes_14_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_13_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_13_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_13_io_to_pes_15_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_13_io_to_pes_15_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_13_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_13_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_13_io_to_pes_16_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_13_io_to_pes_16_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_13_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_13_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_13_io_to_pes_17_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_13_io_to_pes_17_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_13_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_13_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_13_io_to_pes_18_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_13_io_to_pes_18_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_13_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_13_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_13_io_to_pes_19_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_13_io_to_pes_19_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_13_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_13_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_13_io_to_pes_20_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_13_io_to_pes_20_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_13_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_13_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_13_io_to_pes_21_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_13_io_to_pes_21_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_13_io_to_pes_21_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_13_io_to_pes_21_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_13_io_to_pes_22_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_13_io_to_pes_22_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_13_io_to_pes_22_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_13_io_to_pes_22_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_13_io_to_pes_23_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_13_io_to_pes_23_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_13_io_to_pes_23_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_13_io_to_pes_23_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_13_io_to_pes_24_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_13_io_to_pes_24_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_13_io_to_pes_24_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_13_io_to_pes_24_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_13_io_to_pes_25_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_13_io_to_pes_25_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_13_io_to_pes_25_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_13_io_to_pes_25_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_13_io_to_pes_26_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_13_io_to_pes_26_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_13_io_to_pes_26_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_13_io_to_pes_26_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_13_io_to_pes_27_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_13_io_to_pes_27_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_13_io_to_pes_27_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_13_io_to_pes_27_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_13_io_to_pes_28_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_13_io_to_pes_28_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_13_io_to_pes_28_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_13_io_to_pes_28_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_13_io_to_pes_29_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_13_io_to_pes_29_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_13_io_to_mem_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_13_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_14_io_to_pes_0_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_14_io_to_pes_0_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_14_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_14_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_14_io_to_pes_1_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_14_io_to_pes_1_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_14_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_14_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_14_io_to_pes_2_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_14_io_to_pes_2_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_14_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_14_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_14_io_to_pes_3_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_14_io_to_pes_3_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_14_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_14_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_14_io_to_pes_4_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_14_io_to_pes_4_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_14_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_14_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_14_io_to_pes_5_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_14_io_to_pes_5_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_14_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_14_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_14_io_to_pes_6_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_14_io_to_pes_6_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_14_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_14_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_14_io_to_pes_7_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_14_io_to_pes_7_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_14_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_14_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_14_io_to_pes_8_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_14_io_to_pes_8_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_14_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_14_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_14_io_to_pes_9_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_14_io_to_pes_9_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_14_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_14_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_14_io_to_pes_10_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_14_io_to_pes_10_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_14_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_14_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_14_io_to_pes_11_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_14_io_to_pes_11_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_14_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_14_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_14_io_to_pes_12_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_14_io_to_pes_12_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_14_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_14_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_14_io_to_pes_13_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_14_io_to_pes_13_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_14_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_14_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_14_io_to_pes_14_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_14_io_to_pes_14_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_14_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_14_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_14_io_to_pes_15_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_14_io_to_pes_15_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_14_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_14_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_14_io_to_pes_16_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_14_io_to_pes_16_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_14_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_14_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_14_io_to_pes_17_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_14_io_to_pes_17_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_14_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_14_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_14_io_to_pes_18_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_14_io_to_pes_18_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_14_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_14_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_14_io_to_pes_19_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_14_io_to_pes_19_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_14_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_14_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_14_io_to_pes_20_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_14_io_to_pes_20_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_14_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_14_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_14_io_to_pes_21_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_14_io_to_pes_21_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_14_io_to_pes_21_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_14_io_to_pes_21_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_14_io_to_pes_22_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_14_io_to_pes_22_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_14_io_to_pes_22_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_14_io_to_pes_22_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_14_io_to_pes_23_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_14_io_to_pes_23_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_14_io_to_pes_23_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_14_io_to_pes_23_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_14_io_to_pes_24_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_14_io_to_pes_24_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_14_io_to_pes_24_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_14_io_to_pes_24_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_14_io_to_pes_25_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_14_io_to_pes_25_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_14_io_to_pes_25_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_14_io_to_pes_25_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_14_io_to_pes_26_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_14_io_to_pes_26_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_14_io_to_pes_26_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_14_io_to_pes_26_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_14_io_to_pes_27_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_14_io_to_pes_27_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_14_io_to_pes_27_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_14_io_to_pes_27_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_14_io_to_pes_28_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_14_io_to_pes_28_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_14_io_to_pes_28_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_14_io_to_pes_28_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_14_io_to_pes_29_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_14_io_to_pes_29_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_14_io_to_mem_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_14_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_15_io_to_pes_0_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_15_io_to_pes_0_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_15_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_15_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_15_io_to_pes_1_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_15_io_to_pes_1_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_15_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_15_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_15_io_to_pes_2_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_15_io_to_pes_2_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_15_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_15_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_15_io_to_pes_3_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_15_io_to_pes_3_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_15_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_15_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_15_io_to_pes_4_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_15_io_to_pes_4_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_15_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_15_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_15_io_to_pes_5_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_15_io_to_pes_5_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_15_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_15_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_15_io_to_pes_6_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_15_io_to_pes_6_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_15_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_15_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_15_io_to_pes_7_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_15_io_to_pes_7_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_15_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_15_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_15_io_to_pes_8_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_15_io_to_pes_8_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_15_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_15_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_15_io_to_pes_9_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_15_io_to_pes_9_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_15_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_15_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_15_io_to_pes_10_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_15_io_to_pes_10_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_15_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_15_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_15_io_to_pes_11_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_15_io_to_pes_11_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_15_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_15_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_15_io_to_pes_12_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_15_io_to_pes_12_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_15_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_15_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_15_io_to_pes_13_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_15_io_to_pes_13_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_15_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_15_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_15_io_to_pes_14_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_15_io_to_pes_14_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_15_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_15_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_15_io_to_pes_15_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_15_io_to_pes_15_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_15_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_15_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_15_io_to_pes_16_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_15_io_to_pes_16_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_15_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_15_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_15_io_to_pes_17_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_15_io_to_pes_17_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_15_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_15_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_15_io_to_pes_18_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_15_io_to_pes_18_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_15_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_15_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_15_io_to_pes_19_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_15_io_to_pes_19_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_15_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_15_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_15_io_to_pes_20_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_15_io_to_pes_20_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_15_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_15_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_15_io_to_pes_21_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_15_io_to_pes_21_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_15_io_to_pes_21_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_15_io_to_pes_21_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_15_io_to_pes_22_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_15_io_to_pes_22_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_15_io_to_pes_22_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_15_io_to_pes_22_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_15_io_to_pes_23_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_15_io_to_pes_23_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_15_io_to_pes_23_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_15_io_to_pes_23_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_15_io_to_pes_24_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_15_io_to_pes_24_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_15_io_to_pes_24_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_15_io_to_pes_24_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_15_io_to_pes_25_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_15_io_to_pes_25_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_15_io_to_pes_25_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_15_io_to_pes_25_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_15_io_to_pes_26_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_15_io_to_pes_26_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_15_io_to_pes_26_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_15_io_to_pes_26_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_15_io_to_pes_27_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_15_io_to_pes_27_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_15_io_to_pes_27_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_15_io_to_pes_27_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_15_io_to_pes_28_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_15_io_to_pes_28_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_15_io_to_pes_28_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_15_io_to_pes_28_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_15_io_to_pes_29_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_15_io_to_pes_29_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_15_io_to_mem_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_15_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_16_io_to_pes_0_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_16_io_to_pes_0_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_16_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_16_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_16_io_to_pes_1_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_16_io_to_pes_1_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_16_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_16_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_16_io_to_pes_2_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_16_io_to_pes_2_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_16_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_16_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_16_io_to_pes_3_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_16_io_to_pes_3_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_16_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_16_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_16_io_to_pes_4_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_16_io_to_pes_4_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_16_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_16_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_16_io_to_pes_5_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_16_io_to_pes_5_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_16_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_16_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_16_io_to_pes_6_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_16_io_to_pes_6_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_16_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_16_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_16_io_to_pes_7_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_16_io_to_pes_7_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_16_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_16_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_16_io_to_pes_8_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_16_io_to_pes_8_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_16_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_16_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_16_io_to_pes_9_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_16_io_to_pes_9_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_16_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_16_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_16_io_to_pes_10_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_16_io_to_pes_10_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_16_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_16_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_16_io_to_pes_11_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_16_io_to_pes_11_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_16_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_16_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_16_io_to_pes_12_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_16_io_to_pes_12_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_16_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_16_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_16_io_to_pes_13_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_16_io_to_pes_13_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_16_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_16_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_16_io_to_pes_14_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_16_io_to_pes_14_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_16_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_16_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_16_io_to_pes_15_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_16_io_to_pes_15_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_16_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_16_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_16_io_to_pes_16_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_16_io_to_pes_16_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_16_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_16_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_16_io_to_pes_17_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_16_io_to_pes_17_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_16_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_16_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_16_io_to_pes_18_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_16_io_to_pes_18_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_16_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_16_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_16_io_to_pes_19_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_16_io_to_pes_19_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_16_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_16_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_16_io_to_pes_20_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_16_io_to_pes_20_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_16_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_16_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_16_io_to_pes_21_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_16_io_to_pes_21_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_16_io_to_pes_21_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_16_io_to_pes_21_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_16_io_to_pes_22_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_16_io_to_pes_22_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_16_io_to_pes_22_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_16_io_to_pes_22_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_16_io_to_pes_23_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_16_io_to_pes_23_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_16_io_to_pes_23_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_16_io_to_pes_23_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_16_io_to_pes_24_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_16_io_to_pes_24_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_16_io_to_pes_24_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_16_io_to_pes_24_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_16_io_to_pes_25_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_16_io_to_pes_25_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_16_io_to_pes_25_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_16_io_to_pes_25_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_16_io_to_pes_26_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_16_io_to_pes_26_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_16_io_to_pes_26_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_16_io_to_pes_26_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_16_io_to_pes_27_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_16_io_to_pes_27_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_16_io_to_pes_27_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_16_io_to_pes_27_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_16_io_to_pes_28_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_16_io_to_pes_28_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_16_io_to_pes_28_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_16_io_to_pes_28_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_16_io_to_pes_29_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_16_io_to_pes_29_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_16_io_to_mem_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_16_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_17_io_to_pes_0_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_17_io_to_pes_0_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_17_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_17_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_17_io_to_pes_1_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_17_io_to_pes_1_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_17_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_17_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_17_io_to_pes_2_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_17_io_to_pes_2_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_17_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_17_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_17_io_to_pes_3_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_17_io_to_pes_3_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_17_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_17_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_17_io_to_pes_4_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_17_io_to_pes_4_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_17_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_17_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_17_io_to_pes_5_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_17_io_to_pes_5_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_17_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_17_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_17_io_to_pes_6_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_17_io_to_pes_6_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_17_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_17_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_17_io_to_pes_7_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_17_io_to_pes_7_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_17_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_17_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_17_io_to_pes_8_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_17_io_to_pes_8_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_17_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_17_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_17_io_to_pes_9_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_17_io_to_pes_9_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_17_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_17_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_17_io_to_pes_10_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_17_io_to_pes_10_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_17_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_17_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_17_io_to_pes_11_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_17_io_to_pes_11_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_17_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_17_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_17_io_to_pes_12_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_17_io_to_pes_12_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_17_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_17_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_17_io_to_pes_13_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_17_io_to_pes_13_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_17_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_17_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_17_io_to_pes_14_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_17_io_to_pes_14_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_17_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_17_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_17_io_to_pes_15_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_17_io_to_pes_15_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_17_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_17_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_17_io_to_pes_16_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_17_io_to_pes_16_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_17_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_17_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_17_io_to_pes_17_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_17_io_to_pes_17_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_17_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_17_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_17_io_to_pes_18_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_17_io_to_pes_18_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_17_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_17_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_17_io_to_pes_19_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_17_io_to_pes_19_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_17_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_17_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_17_io_to_pes_20_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_17_io_to_pes_20_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_17_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_17_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_17_io_to_pes_21_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_17_io_to_pes_21_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_17_io_to_pes_21_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_17_io_to_pes_21_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_17_io_to_pes_22_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_17_io_to_pes_22_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_17_io_to_pes_22_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_17_io_to_pes_22_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_17_io_to_pes_23_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_17_io_to_pes_23_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_17_io_to_pes_23_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_17_io_to_pes_23_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_17_io_to_pes_24_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_17_io_to_pes_24_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_17_io_to_pes_24_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_17_io_to_pes_24_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_17_io_to_pes_25_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_17_io_to_pes_25_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_17_io_to_pes_25_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_17_io_to_pes_25_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_17_io_to_pes_26_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_17_io_to_pes_26_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_17_io_to_pes_26_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_17_io_to_pes_26_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_17_io_to_pes_27_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_17_io_to_pes_27_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_17_io_to_pes_27_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_17_io_to_pes_27_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_17_io_to_pes_28_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_17_io_to_pes_28_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_17_io_to_pes_28_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_17_io_to_pes_28_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_17_io_to_pes_29_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_17_io_to_pes_29_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_17_io_to_mem_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_17_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_18_io_to_pes_0_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_18_io_to_pes_0_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_18_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_18_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_18_io_to_pes_1_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_18_io_to_pes_1_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_18_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_18_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_18_io_to_pes_2_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_18_io_to_pes_2_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_18_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_18_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_18_io_to_pes_3_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_18_io_to_pes_3_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_18_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_18_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_18_io_to_pes_4_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_18_io_to_pes_4_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_18_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_18_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_18_io_to_pes_5_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_18_io_to_pes_5_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_18_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_18_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_18_io_to_pes_6_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_18_io_to_pes_6_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_18_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_18_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_18_io_to_pes_7_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_18_io_to_pes_7_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_18_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_18_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_18_io_to_pes_8_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_18_io_to_pes_8_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_18_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_18_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_18_io_to_pes_9_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_18_io_to_pes_9_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_18_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_18_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_18_io_to_pes_10_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_18_io_to_pes_10_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_18_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_18_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_18_io_to_pes_11_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_18_io_to_pes_11_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_18_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_18_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_18_io_to_pes_12_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_18_io_to_pes_12_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_18_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_18_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_18_io_to_pes_13_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_18_io_to_pes_13_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_18_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_18_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_18_io_to_pes_14_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_18_io_to_pes_14_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_18_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_18_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_18_io_to_pes_15_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_18_io_to_pes_15_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_18_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_18_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_18_io_to_pes_16_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_18_io_to_pes_16_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_18_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_18_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_18_io_to_pes_17_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_18_io_to_pes_17_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_18_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_18_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_18_io_to_pes_18_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_18_io_to_pes_18_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_18_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_18_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_18_io_to_pes_19_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_18_io_to_pes_19_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_18_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_18_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_18_io_to_pes_20_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_18_io_to_pes_20_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_18_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_18_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_18_io_to_pes_21_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_18_io_to_pes_21_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_18_io_to_pes_21_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_18_io_to_pes_21_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_18_io_to_pes_22_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_18_io_to_pes_22_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_18_io_to_pes_22_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_18_io_to_pes_22_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_18_io_to_pes_23_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_18_io_to_pes_23_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_18_io_to_pes_23_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_18_io_to_pes_23_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_18_io_to_pes_24_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_18_io_to_pes_24_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_18_io_to_pes_24_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_18_io_to_pes_24_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_18_io_to_pes_25_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_18_io_to_pes_25_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_18_io_to_pes_25_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_18_io_to_pes_25_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_18_io_to_pes_26_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_18_io_to_pes_26_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_18_io_to_pes_26_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_18_io_to_pes_26_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_18_io_to_pes_27_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_18_io_to_pes_27_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_18_io_to_pes_27_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_18_io_to_pes_27_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_18_io_to_pes_28_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_18_io_to_pes_28_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_18_io_to_pes_28_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_18_io_to_pes_28_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_18_io_to_pes_29_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_18_io_to_pes_29_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_18_io_to_mem_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_18_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_19_io_to_pes_0_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_19_io_to_pes_0_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_19_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_19_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_19_io_to_pes_1_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_19_io_to_pes_1_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_19_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_19_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_19_io_to_pes_2_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_19_io_to_pes_2_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_19_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_19_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_19_io_to_pes_3_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_19_io_to_pes_3_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_19_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_19_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_19_io_to_pes_4_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_19_io_to_pes_4_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_19_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_19_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_19_io_to_pes_5_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_19_io_to_pes_5_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_19_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_19_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_19_io_to_pes_6_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_19_io_to_pes_6_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_19_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_19_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_19_io_to_pes_7_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_19_io_to_pes_7_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_19_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_19_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_19_io_to_pes_8_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_19_io_to_pes_8_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_19_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_19_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_19_io_to_pes_9_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_19_io_to_pes_9_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_19_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_19_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_19_io_to_pes_10_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_19_io_to_pes_10_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_19_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_19_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_19_io_to_pes_11_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_19_io_to_pes_11_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_19_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_19_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_19_io_to_pes_12_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_19_io_to_pes_12_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_19_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_19_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_19_io_to_pes_13_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_19_io_to_pes_13_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_19_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_19_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_19_io_to_pes_14_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_19_io_to_pes_14_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_19_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_19_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_19_io_to_pes_15_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_19_io_to_pes_15_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_19_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_19_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_19_io_to_pes_16_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_19_io_to_pes_16_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_19_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_19_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_19_io_to_pes_17_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_19_io_to_pes_17_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_19_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_19_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_19_io_to_pes_18_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_19_io_to_pes_18_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_19_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_19_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_19_io_to_pes_19_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_19_io_to_pes_19_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_19_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_19_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_19_io_to_pes_20_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_19_io_to_pes_20_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_19_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_19_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_19_io_to_pes_21_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_19_io_to_pes_21_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_19_io_to_pes_21_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_19_io_to_pes_21_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_19_io_to_pes_22_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_19_io_to_pes_22_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_19_io_to_pes_22_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_19_io_to_pes_22_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_19_io_to_pes_23_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_19_io_to_pes_23_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_19_io_to_pes_23_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_19_io_to_pes_23_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_19_io_to_pes_24_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_19_io_to_pes_24_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_19_io_to_pes_24_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_19_io_to_pes_24_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_19_io_to_pes_25_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_19_io_to_pes_25_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_19_io_to_pes_25_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_19_io_to_pes_25_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_19_io_to_pes_26_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_19_io_to_pes_26_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_19_io_to_pes_26_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_19_io_to_pes_26_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_19_io_to_pes_27_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_19_io_to_pes_27_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_19_io_to_pes_27_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_19_io_to_pes_27_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_19_io_to_pes_28_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_19_io_to_pes_28_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_19_io_to_pes_28_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_19_io_to_pes_28_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_19_io_to_pes_29_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_19_io_to_pes_29_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_19_io_to_mem_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_19_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_20_io_to_pes_0_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_20_io_to_pes_0_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_20_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_20_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_20_io_to_pes_1_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_20_io_to_pes_1_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_20_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_20_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_20_io_to_pes_2_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_20_io_to_pes_2_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_20_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_20_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_20_io_to_pes_3_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_20_io_to_pes_3_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_20_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_20_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_20_io_to_pes_4_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_20_io_to_pes_4_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_20_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_20_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_20_io_to_pes_5_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_20_io_to_pes_5_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_20_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_20_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_20_io_to_pes_6_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_20_io_to_pes_6_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_20_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_20_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_20_io_to_pes_7_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_20_io_to_pes_7_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_20_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_20_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_20_io_to_pes_8_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_20_io_to_pes_8_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_20_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_20_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_20_io_to_pes_9_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_20_io_to_pes_9_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_20_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_20_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_20_io_to_pes_10_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_20_io_to_pes_10_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_20_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_20_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_20_io_to_pes_11_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_20_io_to_pes_11_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_20_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_20_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_20_io_to_pes_12_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_20_io_to_pes_12_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_20_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_20_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_20_io_to_pes_13_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_20_io_to_pes_13_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_20_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_20_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_20_io_to_pes_14_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_20_io_to_pes_14_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_20_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_20_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_20_io_to_pes_15_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_20_io_to_pes_15_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_20_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_20_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_20_io_to_pes_16_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_20_io_to_pes_16_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_20_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_20_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_20_io_to_pes_17_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_20_io_to_pes_17_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_20_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_20_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_20_io_to_pes_18_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_20_io_to_pes_18_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_20_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_20_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_20_io_to_pes_19_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_20_io_to_pes_19_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_20_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_20_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_20_io_to_pes_20_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_20_io_to_pes_20_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_20_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_20_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_20_io_to_pes_21_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_20_io_to_pes_21_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_20_io_to_pes_21_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_20_io_to_pes_21_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_20_io_to_pes_22_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_20_io_to_pes_22_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_20_io_to_pes_22_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_20_io_to_pes_22_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_20_io_to_pes_23_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_20_io_to_pes_23_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_20_io_to_pes_23_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_20_io_to_pes_23_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_20_io_to_pes_24_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_20_io_to_pes_24_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_20_io_to_pes_24_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_20_io_to_pes_24_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_20_io_to_pes_25_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_20_io_to_pes_25_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_20_io_to_pes_25_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_20_io_to_pes_25_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_20_io_to_pes_26_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_20_io_to_pes_26_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_20_io_to_pes_26_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_20_io_to_pes_26_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_20_io_to_pes_27_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_20_io_to_pes_27_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_20_io_to_pes_27_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_20_io_to_pes_27_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_20_io_to_pes_28_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_20_io_to_pes_28_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_20_io_to_pes_28_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_20_io_to_pes_28_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_20_io_to_pes_29_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_20_io_to_pes_29_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_20_io_to_mem_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_20_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_21_io_to_pes_0_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_21_io_to_pes_0_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_21_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_21_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_21_io_to_pes_1_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_21_io_to_pes_1_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_21_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_21_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_21_io_to_pes_2_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_21_io_to_pes_2_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_21_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_21_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_21_io_to_pes_3_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_21_io_to_pes_3_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_21_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_21_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_21_io_to_pes_4_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_21_io_to_pes_4_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_21_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_21_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_21_io_to_pes_5_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_21_io_to_pes_5_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_21_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_21_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_21_io_to_pes_6_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_21_io_to_pes_6_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_21_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_21_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_21_io_to_pes_7_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_21_io_to_pes_7_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_21_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_21_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_21_io_to_pes_8_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_21_io_to_pes_8_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_21_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_21_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_21_io_to_pes_9_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_21_io_to_pes_9_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_21_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_21_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_21_io_to_pes_10_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_21_io_to_pes_10_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_21_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_21_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_21_io_to_pes_11_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_21_io_to_pes_11_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_21_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_21_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_21_io_to_pes_12_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_21_io_to_pes_12_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_21_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_21_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_21_io_to_pes_13_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_21_io_to_pes_13_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_21_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_21_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_21_io_to_pes_14_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_21_io_to_pes_14_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_21_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_21_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_21_io_to_pes_15_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_21_io_to_pes_15_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_21_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_21_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_21_io_to_pes_16_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_21_io_to_pes_16_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_21_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_21_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_21_io_to_pes_17_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_21_io_to_pes_17_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_21_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_21_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_21_io_to_pes_18_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_21_io_to_pes_18_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_21_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_21_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_21_io_to_pes_19_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_21_io_to_pes_19_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_21_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_21_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_21_io_to_pes_20_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_21_io_to_pes_20_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_21_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_21_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_21_io_to_pes_21_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_21_io_to_pes_21_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_21_io_to_pes_21_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_21_io_to_pes_21_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_21_io_to_pes_22_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_21_io_to_pes_22_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_21_io_to_pes_22_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_21_io_to_pes_22_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_21_io_to_pes_23_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_21_io_to_pes_23_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_21_io_to_pes_23_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_21_io_to_pes_23_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_21_io_to_pes_24_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_21_io_to_pes_24_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_21_io_to_pes_24_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_21_io_to_pes_24_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_21_io_to_pes_25_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_21_io_to_pes_25_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_21_io_to_pes_25_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_21_io_to_pes_25_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_21_io_to_pes_26_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_21_io_to_pes_26_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_21_io_to_pes_26_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_21_io_to_pes_26_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_21_io_to_pes_27_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_21_io_to_pes_27_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_21_io_to_pes_27_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_21_io_to_pes_27_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_21_io_to_pes_28_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_21_io_to_pes_28_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_21_io_to_pes_28_out_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_21_io_to_pes_28_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_21_io_to_pes_29_in_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_21_io_to_pes_29_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_21_io_to_mem_valid; // @[pe.scala 229:13]
  wire [15:0] PENetwork_21_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_22_io_to_pes_0_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_22_io_to_pes_0_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_22_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_22_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_22_io_to_pes_1_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_22_io_to_pes_1_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_22_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_22_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_22_io_to_pes_2_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_22_io_to_pes_2_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_22_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_22_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_22_io_to_pes_3_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_22_io_to_pes_3_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_22_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_22_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_22_io_to_pes_4_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_22_io_to_pes_4_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_22_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_22_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_22_io_to_pes_5_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_22_io_to_pes_5_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_22_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_22_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_22_io_to_pes_6_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_22_io_to_pes_6_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_22_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_22_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_22_io_to_pes_7_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_22_io_to_pes_7_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_22_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_22_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_22_io_to_pes_8_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_22_io_to_pes_8_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_22_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_22_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_22_io_to_pes_9_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_22_io_to_pes_9_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_22_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_22_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_22_io_to_pes_10_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_22_io_to_pes_10_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_22_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_22_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_22_io_to_pes_11_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_22_io_to_pes_11_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_22_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_22_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_22_io_to_pes_12_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_22_io_to_pes_12_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_22_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_22_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_22_io_to_pes_13_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_22_io_to_pes_13_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_22_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_22_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_22_io_to_pes_14_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_22_io_to_pes_14_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_22_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_22_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_22_io_to_pes_15_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_22_io_to_pes_15_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_22_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_22_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_22_io_to_pes_16_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_22_io_to_pes_16_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_22_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_22_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_22_io_to_pes_17_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_22_io_to_pes_17_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_22_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_22_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_22_io_to_pes_18_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_22_io_to_pes_18_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_22_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_22_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_22_io_to_pes_19_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_22_io_to_pes_19_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_22_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_22_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_22_io_to_pes_20_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_22_io_to_pes_20_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_22_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_22_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_22_io_to_pes_21_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_22_io_to_pes_21_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_22_io_to_mem_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_22_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_23_io_to_pes_0_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_23_io_to_pes_0_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_23_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_23_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_23_io_to_pes_1_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_23_io_to_pes_1_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_23_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_23_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_23_io_to_pes_2_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_23_io_to_pes_2_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_23_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_23_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_23_io_to_pes_3_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_23_io_to_pes_3_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_23_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_23_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_23_io_to_pes_4_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_23_io_to_pes_4_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_23_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_23_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_23_io_to_pes_5_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_23_io_to_pes_5_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_23_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_23_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_23_io_to_pes_6_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_23_io_to_pes_6_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_23_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_23_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_23_io_to_pes_7_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_23_io_to_pes_7_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_23_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_23_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_23_io_to_pes_8_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_23_io_to_pes_8_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_23_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_23_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_23_io_to_pes_9_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_23_io_to_pes_9_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_23_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_23_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_23_io_to_pes_10_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_23_io_to_pes_10_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_23_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_23_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_23_io_to_pes_11_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_23_io_to_pes_11_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_23_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_23_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_23_io_to_pes_12_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_23_io_to_pes_12_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_23_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_23_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_23_io_to_pes_13_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_23_io_to_pes_13_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_23_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_23_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_23_io_to_pes_14_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_23_io_to_pes_14_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_23_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_23_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_23_io_to_pes_15_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_23_io_to_pes_15_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_23_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_23_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_23_io_to_pes_16_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_23_io_to_pes_16_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_23_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_23_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_23_io_to_pes_17_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_23_io_to_pes_17_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_23_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_23_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_23_io_to_pes_18_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_23_io_to_pes_18_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_23_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_23_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_23_io_to_pes_19_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_23_io_to_pes_19_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_23_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_23_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_23_io_to_pes_20_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_23_io_to_pes_20_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_23_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_23_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_23_io_to_pes_21_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_23_io_to_pes_21_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_23_io_to_mem_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_23_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_24_io_to_pes_0_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_24_io_to_pes_0_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_24_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_24_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_24_io_to_pes_1_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_24_io_to_pes_1_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_24_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_24_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_24_io_to_pes_2_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_24_io_to_pes_2_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_24_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_24_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_24_io_to_pes_3_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_24_io_to_pes_3_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_24_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_24_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_24_io_to_pes_4_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_24_io_to_pes_4_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_24_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_24_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_24_io_to_pes_5_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_24_io_to_pes_5_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_24_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_24_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_24_io_to_pes_6_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_24_io_to_pes_6_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_24_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_24_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_24_io_to_pes_7_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_24_io_to_pes_7_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_24_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_24_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_24_io_to_pes_8_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_24_io_to_pes_8_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_24_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_24_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_24_io_to_pes_9_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_24_io_to_pes_9_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_24_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_24_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_24_io_to_pes_10_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_24_io_to_pes_10_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_24_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_24_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_24_io_to_pes_11_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_24_io_to_pes_11_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_24_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_24_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_24_io_to_pes_12_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_24_io_to_pes_12_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_24_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_24_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_24_io_to_pes_13_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_24_io_to_pes_13_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_24_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_24_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_24_io_to_pes_14_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_24_io_to_pes_14_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_24_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_24_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_24_io_to_pes_15_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_24_io_to_pes_15_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_24_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_24_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_24_io_to_pes_16_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_24_io_to_pes_16_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_24_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_24_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_24_io_to_pes_17_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_24_io_to_pes_17_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_24_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_24_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_24_io_to_pes_18_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_24_io_to_pes_18_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_24_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_24_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_24_io_to_pes_19_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_24_io_to_pes_19_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_24_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_24_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_24_io_to_pes_20_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_24_io_to_pes_20_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_24_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_24_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_24_io_to_pes_21_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_24_io_to_pes_21_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_24_io_to_mem_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_24_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_25_io_to_pes_0_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_25_io_to_pes_0_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_25_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_25_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_25_io_to_pes_1_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_25_io_to_pes_1_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_25_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_25_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_25_io_to_pes_2_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_25_io_to_pes_2_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_25_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_25_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_25_io_to_pes_3_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_25_io_to_pes_3_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_25_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_25_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_25_io_to_pes_4_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_25_io_to_pes_4_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_25_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_25_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_25_io_to_pes_5_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_25_io_to_pes_5_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_25_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_25_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_25_io_to_pes_6_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_25_io_to_pes_6_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_25_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_25_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_25_io_to_pes_7_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_25_io_to_pes_7_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_25_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_25_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_25_io_to_pes_8_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_25_io_to_pes_8_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_25_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_25_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_25_io_to_pes_9_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_25_io_to_pes_9_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_25_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_25_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_25_io_to_pes_10_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_25_io_to_pes_10_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_25_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_25_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_25_io_to_pes_11_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_25_io_to_pes_11_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_25_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_25_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_25_io_to_pes_12_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_25_io_to_pes_12_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_25_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_25_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_25_io_to_pes_13_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_25_io_to_pes_13_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_25_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_25_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_25_io_to_pes_14_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_25_io_to_pes_14_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_25_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_25_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_25_io_to_pes_15_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_25_io_to_pes_15_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_25_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_25_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_25_io_to_pes_16_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_25_io_to_pes_16_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_25_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_25_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_25_io_to_pes_17_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_25_io_to_pes_17_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_25_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_25_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_25_io_to_pes_18_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_25_io_to_pes_18_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_25_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_25_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_25_io_to_pes_19_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_25_io_to_pes_19_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_25_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_25_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_25_io_to_pes_20_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_25_io_to_pes_20_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_25_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_25_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_25_io_to_pes_21_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_25_io_to_pes_21_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_25_io_to_mem_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_25_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_26_io_to_pes_0_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_26_io_to_pes_0_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_26_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_26_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_26_io_to_pes_1_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_26_io_to_pes_1_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_26_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_26_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_26_io_to_pes_2_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_26_io_to_pes_2_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_26_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_26_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_26_io_to_pes_3_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_26_io_to_pes_3_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_26_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_26_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_26_io_to_pes_4_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_26_io_to_pes_4_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_26_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_26_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_26_io_to_pes_5_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_26_io_to_pes_5_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_26_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_26_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_26_io_to_pes_6_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_26_io_to_pes_6_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_26_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_26_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_26_io_to_pes_7_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_26_io_to_pes_7_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_26_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_26_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_26_io_to_pes_8_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_26_io_to_pes_8_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_26_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_26_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_26_io_to_pes_9_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_26_io_to_pes_9_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_26_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_26_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_26_io_to_pes_10_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_26_io_to_pes_10_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_26_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_26_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_26_io_to_pes_11_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_26_io_to_pes_11_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_26_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_26_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_26_io_to_pes_12_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_26_io_to_pes_12_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_26_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_26_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_26_io_to_pes_13_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_26_io_to_pes_13_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_26_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_26_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_26_io_to_pes_14_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_26_io_to_pes_14_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_26_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_26_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_26_io_to_pes_15_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_26_io_to_pes_15_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_26_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_26_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_26_io_to_pes_16_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_26_io_to_pes_16_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_26_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_26_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_26_io_to_pes_17_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_26_io_to_pes_17_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_26_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_26_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_26_io_to_pes_18_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_26_io_to_pes_18_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_26_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_26_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_26_io_to_pes_19_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_26_io_to_pes_19_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_26_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_26_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_26_io_to_pes_20_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_26_io_to_pes_20_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_26_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_26_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_26_io_to_pes_21_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_26_io_to_pes_21_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_26_io_to_mem_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_26_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_27_io_to_pes_0_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_27_io_to_pes_0_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_27_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_27_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_27_io_to_pes_1_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_27_io_to_pes_1_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_27_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_27_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_27_io_to_pes_2_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_27_io_to_pes_2_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_27_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_27_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_27_io_to_pes_3_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_27_io_to_pes_3_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_27_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_27_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_27_io_to_pes_4_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_27_io_to_pes_4_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_27_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_27_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_27_io_to_pes_5_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_27_io_to_pes_5_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_27_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_27_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_27_io_to_pes_6_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_27_io_to_pes_6_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_27_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_27_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_27_io_to_pes_7_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_27_io_to_pes_7_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_27_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_27_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_27_io_to_pes_8_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_27_io_to_pes_8_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_27_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_27_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_27_io_to_pes_9_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_27_io_to_pes_9_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_27_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_27_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_27_io_to_pes_10_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_27_io_to_pes_10_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_27_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_27_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_27_io_to_pes_11_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_27_io_to_pes_11_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_27_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_27_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_27_io_to_pes_12_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_27_io_to_pes_12_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_27_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_27_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_27_io_to_pes_13_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_27_io_to_pes_13_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_27_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_27_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_27_io_to_pes_14_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_27_io_to_pes_14_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_27_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_27_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_27_io_to_pes_15_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_27_io_to_pes_15_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_27_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_27_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_27_io_to_pes_16_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_27_io_to_pes_16_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_27_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_27_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_27_io_to_pes_17_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_27_io_to_pes_17_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_27_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_27_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_27_io_to_pes_18_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_27_io_to_pes_18_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_27_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_27_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_27_io_to_pes_19_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_27_io_to_pes_19_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_27_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_27_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_27_io_to_pes_20_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_27_io_to_pes_20_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_27_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_27_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_27_io_to_pes_21_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_27_io_to_pes_21_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_27_io_to_mem_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_27_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_28_io_to_pes_0_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_28_io_to_pes_0_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_28_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_28_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_28_io_to_pes_1_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_28_io_to_pes_1_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_28_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_28_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_28_io_to_pes_2_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_28_io_to_pes_2_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_28_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_28_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_28_io_to_pes_3_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_28_io_to_pes_3_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_28_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_28_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_28_io_to_pes_4_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_28_io_to_pes_4_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_28_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_28_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_28_io_to_pes_5_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_28_io_to_pes_5_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_28_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_28_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_28_io_to_pes_6_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_28_io_to_pes_6_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_28_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_28_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_28_io_to_pes_7_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_28_io_to_pes_7_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_28_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_28_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_28_io_to_pes_8_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_28_io_to_pes_8_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_28_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_28_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_28_io_to_pes_9_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_28_io_to_pes_9_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_28_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_28_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_28_io_to_pes_10_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_28_io_to_pes_10_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_28_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_28_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_28_io_to_pes_11_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_28_io_to_pes_11_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_28_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_28_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_28_io_to_pes_12_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_28_io_to_pes_12_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_28_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_28_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_28_io_to_pes_13_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_28_io_to_pes_13_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_28_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_28_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_28_io_to_pes_14_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_28_io_to_pes_14_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_28_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_28_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_28_io_to_pes_15_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_28_io_to_pes_15_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_28_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_28_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_28_io_to_pes_16_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_28_io_to_pes_16_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_28_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_28_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_28_io_to_pes_17_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_28_io_to_pes_17_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_28_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_28_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_28_io_to_pes_18_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_28_io_to_pes_18_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_28_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_28_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_28_io_to_pes_19_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_28_io_to_pes_19_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_28_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_28_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_28_io_to_pes_20_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_28_io_to_pes_20_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_28_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_28_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_28_io_to_pes_21_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_28_io_to_pes_21_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_28_io_to_mem_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_28_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_29_io_to_pes_0_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_29_io_to_pes_0_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_29_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_29_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_29_io_to_pes_1_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_29_io_to_pes_1_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_29_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_29_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_29_io_to_pes_2_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_29_io_to_pes_2_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_29_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_29_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_29_io_to_pes_3_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_29_io_to_pes_3_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_29_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_29_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_29_io_to_pes_4_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_29_io_to_pes_4_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_29_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_29_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_29_io_to_pes_5_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_29_io_to_pes_5_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_29_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_29_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_29_io_to_pes_6_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_29_io_to_pes_6_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_29_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_29_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_29_io_to_pes_7_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_29_io_to_pes_7_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_29_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_29_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_29_io_to_pes_8_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_29_io_to_pes_8_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_29_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_29_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_29_io_to_pes_9_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_29_io_to_pes_9_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_29_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_29_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_29_io_to_pes_10_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_29_io_to_pes_10_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_29_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_29_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_29_io_to_pes_11_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_29_io_to_pes_11_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_29_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_29_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_29_io_to_pes_12_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_29_io_to_pes_12_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_29_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_29_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_29_io_to_pes_13_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_29_io_to_pes_13_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_29_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_29_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_29_io_to_pes_14_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_29_io_to_pes_14_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_29_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_29_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_29_io_to_pes_15_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_29_io_to_pes_15_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_29_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_29_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_29_io_to_pes_16_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_29_io_to_pes_16_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_29_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_29_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_29_io_to_pes_17_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_29_io_to_pes_17_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_29_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_29_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_29_io_to_pes_18_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_29_io_to_pes_18_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_29_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_29_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_29_io_to_pes_19_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_29_io_to_pes_19_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_29_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_29_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_29_io_to_pes_20_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_29_io_to_pes_20_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_29_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_29_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_29_io_to_pes_21_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_29_io_to_pes_21_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_29_io_to_mem_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_29_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_30_io_to_pes_0_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_30_io_to_pes_0_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_30_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_30_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_30_io_to_pes_1_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_30_io_to_pes_1_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_30_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_30_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_30_io_to_pes_2_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_30_io_to_pes_2_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_30_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_30_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_30_io_to_pes_3_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_30_io_to_pes_3_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_30_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_30_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_30_io_to_pes_4_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_30_io_to_pes_4_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_30_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_30_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_30_io_to_pes_5_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_30_io_to_pes_5_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_30_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_30_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_30_io_to_pes_6_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_30_io_to_pes_6_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_30_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_30_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_30_io_to_pes_7_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_30_io_to_pes_7_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_30_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_30_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_30_io_to_pes_8_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_30_io_to_pes_8_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_30_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_30_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_30_io_to_pes_9_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_30_io_to_pes_9_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_30_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_30_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_30_io_to_pes_10_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_30_io_to_pes_10_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_30_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_30_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_30_io_to_pes_11_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_30_io_to_pes_11_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_30_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_30_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_30_io_to_pes_12_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_30_io_to_pes_12_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_30_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_30_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_30_io_to_pes_13_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_30_io_to_pes_13_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_30_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_30_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_30_io_to_pes_14_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_30_io_to_pes_14_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_30_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_30_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_30_io_to_pes_15_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_30_io_to_pes_15_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_30_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_30_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_30_io_to_pes_16_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_30_io_to_pes_16_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_30_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_30_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_30_io_to_pes_17_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_30_io_to_pes_17_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_30_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_30_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_30_io_to_pes_18_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_30_io_to_pes_18_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_30_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_30_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_30_io_to_pes_19_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_30_io_to_pes_19_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_30_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_30_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_30_io_to_pes_20_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_30_io_to_pes_20_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_30_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_30_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_30_io_to_pes_21_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_30_io_to_pes_21_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_30_io_to_mem_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_30_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_31_io_to_pes_0_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_31_io_to_pes_0_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_31_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_31_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_31_io_to_pes_1_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_31_io_to_pes_1_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_31_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_31_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_31_io_to_pes_2_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_31_io_to_pes_2_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_31_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_31_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_31_io_to_pes_3_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_31_io_to_pes_3_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_31_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_31_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_31_io_to_pes_4_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_31_io_to_pes_4_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_31_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_31_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_31_io_to_pes_5_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_31_io_to_pes_5_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_31_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_31_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_31_io_to_pes_6_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_31_io_to_pes_6_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_31_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_31_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_31_io_to_pes_7_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_31_io_to_pes_7_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_31_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_31_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_31_io_to_pes_8_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_31_io_to_pes_8_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_31_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_31_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_31_io_to_pes_9_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_31_io_to_pes_9_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_31_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_31_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_31_io_to_pes_10_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_31_io_to_pes_10_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_31_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_31_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_31_io_to_pes_11_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_31_io_to_pes_11_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_31_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_31_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_31_io_to_pes_12_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_31_io_to_pes_12_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_31_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_31_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_31_io_to_pes_13_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_31_io_to_pes_13_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_31_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_31_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_31_io_to_pes_14_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_31_io_to_pes_14_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_31_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_31_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_31_io_to_pes_15_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_31_io_to_pes_15_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_31_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_31_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_31_io_to_pes_16_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_31_io_to_pes_16_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_31_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_31_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_31_io_to_pes_17_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_31_io_to_pes_17_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_31_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_31_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_31_io_to_pes_18_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_31_io_to_pes_18_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_31_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_31_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_31_io_to_pes_19_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_31_io_to_pes_19_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_31_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_31_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_31_io_to_pes_20_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_31_io_to_pes_20_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_31_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_31_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_31_io_to_pes_21_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_31_io_to_pes_21_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_31_io_to_mem_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_31_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_32_io_to_pes_0_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_32_io_to_pes_0_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_32_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_32_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_32_io_to_pes_1_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_32_io_to_pes_1_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_32_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_32_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_32_io_to_pes_2_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_32_io_to_pes_2_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_32_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_32_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_32_io_to_pes_3_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_32_io_to_pes_3_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_32_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_32_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_32_io_to_pes_4_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_32_io_to_pes_4_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_32_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_32_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_32_io_to_pes_5_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_32_io_to_pes_5_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_32_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_32_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_32_io_to_pes_6_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_32_io_to_pes_6_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_32_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_32_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_32_io_to_pes_7_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_32_io_to_pes_7_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_32_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_32_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_32_io_to_pes_8_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_32_io_to_pes_8_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_32_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_32_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_32_io_to_pes_9_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_32_io_to_pes_9_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_32_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_32_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_32_io_to_pes_10_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_32_io_to_pes_10_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_32_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_32_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_32_io_to_pes_11_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_32_io_to_pes_11_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_32_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_32_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_32_io_to_pes_12_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_32_io_to_pes_12_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_32_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_32_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_32_io_to_pes_13_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_32_io_to_pes_13_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_32_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_32_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_32_io_to_pes_14_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_32_io_to_pes_14_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_32_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_32_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_32_io_to_pes_15_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_32_io_to_pes_15_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_32_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_32_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_32_io_to_pes_16_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_32_io_to_pes_16_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_32_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_32_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_32_io_to_pes_17_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_32_io_to_pes_17_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_32_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_32_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_32_io_to_pes_18_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_32_io_to_pes_18_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_32_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_32_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_32_io_to_pes_19_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_32_io_to_pes_19_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_32_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_32_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_32_io_to_pes_20_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_32_io_to_pes_20_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_32_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_32_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_32_io_to_pes_21_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_32_io_to_pes_21_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_32_io_to_mem_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_32_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_33_io_to_pes_0_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_33_io_to_pes_0_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_33_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_33_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_33_io_to_pes_1_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_33_io_to_pes_1_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_33_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_33_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_33_io_to_pes_2_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_33_io_to_pes_2_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_33_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_33_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_33_io_to_pes_3_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_33_io_to_pes_3_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_33_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_33_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_33_io_to_pes_4_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_33_io_to_pes_4_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_33_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_33_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_33_io_to_pes_5_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_33_io_to_pes_5_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_33_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_33_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_33_io_to_pes_6_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_33_io_to_pes_6_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_33_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_33_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_33_io_to_pes_7_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_33_io_to_pes_7_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_33_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_33_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_33_io_to_pes_8_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_33_io_to_pes_8_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_33_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_33_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_33_io_to_pes_9_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_33_io_to_pes_9_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_33_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_33_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_33_io_to_pes_10_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_33_io_to_pes_10_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_33_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_33_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_33_io_to_pes_11_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_33_io_to_pes_11_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_33_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_33_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_33_io_to_pes_12_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_33_io_to_pes_12_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_33_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_33_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_33_io_to_pes_13_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_33_io_to_pes_13_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_33_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_33_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_33_io_to_pes_14_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_33_io_to_pes_14_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_33_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_33_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_33_io_to_pes_15_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_33_io_to_pes_15_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_33_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_33_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_33_io_to_pes_16_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_33_io_to_pes_16_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_33_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_33_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_33_io_to_pes_17_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_33_io_to_pes_17_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_33_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_33_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_33_io_to_pes_18_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_33_io_to_pes_18_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_33_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_33_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_33_io_to_pes_19_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_33_io_to_pes_19_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_33_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_33_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_33_io_to_pes_20_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_33_io_to_pes_20_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_33_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_33_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_33_io_to_pes_21_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_33_io_to_pes_21_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_33_io_to_mem_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_33_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_34_io_to_pes_0_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_34_io_to_pes_0_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_34_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_34_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_34_io_to_pes_1_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_34_io_to_pes_1_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_34_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_34_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_34_io_to_pes_2_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_34_io_to_pes_2_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_34_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_34_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_34_io_to_pes_3_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_34_io_to_pes_3_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_34_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_34_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_34_io_to_pes_4_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_34_io_to_pes_4_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_34_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_34_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_34_io_to_pes_5_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_34_io_to_pes_5_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_34_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_34_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_34_io_to_pes_6_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_34_io_to_pes_6_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_34_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_34_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_34_io_to_pes_7_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_34_io_to_pes_7_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_34_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_34_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_34_io_to_pes_8_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_34_io_to_pes_8_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_34_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_34_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_34_io_to_pes_9_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_34_io_to_pes_9_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_34_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_34_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_34_io_to_pes_10_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_34_io_to_pes_10_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_34_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_34_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_34_io_to_pes_11_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_34_io_to_pes_11_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_34_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_34_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_34_io_to_pes_12_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_34_io_to_pes_12_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_34_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_34_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_34_io_to_pes_13_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_34_io_to_pes_13_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_34_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_34_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_34_io_to_pes_14_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_34_io_to_pes_14_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_34_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_34_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_34_io_to_pes_15_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_34_io_to_pes_15_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_34_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_34_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_34_io_to_pes_16_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_34_io_to_pes_16_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_34_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_34_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_34_io_to_pes_17_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_34_io_to_pes_17_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_34_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_34_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_34_io_to_pes_18_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_34_io_to_pes_18_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_34_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_34_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_34_io_to_pes_19_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_34_io_to_pes_19_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_34_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_34_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_34_io_to_pes_20_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_34_io_to_pes_20_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_34_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_34_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_34_io_to_pes_21_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_34_io_to_pes_21_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_34_io_to_mem_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_34_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_35_io_to_pes_0_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_35_io_to_pes_0_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_35_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_35_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_35_io_to_pes_1_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_35_io_to_pes_1_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_35_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_35_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_35_io_to_pes_2_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_35_io_to_pes_2_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_35_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_35_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_35_io_to_pes_3_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_35_io_to_pes_3_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_35_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_35_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_35_io_to_pes_4_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_35_io_to_pes_4_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_35_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_35_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_35_io_to_pes_5_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_35_io_to_pes_5_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_35_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_35_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_35_io_to_pes_6_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_35_io_to_pes_6_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_35_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_35_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_35_io_to_pes_7_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_35_io_to_pes_7_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_35_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_35_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_35_io_to_pes_8_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_35_io_to_pes_8_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_35_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_35_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_35_io_to_pes_9_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_35_io_to_pes_9_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_35_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_35_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_35_io_to_pes_10_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_35_io_to_pes_10_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_35_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_35_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_35_io_to_pes_11_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_35_io_to_pes_11_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_35_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_35_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_35_io_to_pes_12_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_35_io_to_pes_12_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_35_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_35_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_35_io_to_pes_13_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_35_io_to_pes_13_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_35_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_35_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_35_io_to_pes_14_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_35_io_to_pes_14_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_35_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_35_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_35_io_to_pes_15_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_35_io_to_pes_15_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_35_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_35_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_35_io_to_pes_16_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_35_io_to_pes_16_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_35_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_35_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_35_io_to_pes_17_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_35_io_to_pes_17_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_35_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_35_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_35_io_to_pes_18_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_35_io_to_pes_18_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_35_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_35_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_35_io_to_pes_19_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_35_io_to_pes_19_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_35_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_35_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_35_io_to_pes_20_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_35_io_to_pes_20_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_35_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_35_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_35_io_to_pes_21_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_35_io_to_pes_21_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_35_io_to_mem_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_35_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_36_io_to_pes_0_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_36_io_to_pes_0_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_36_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_36_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_36_io_to_pes_1_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_36_io_to_pes_1_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_36_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_36_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_36_io_to_pes_2_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_36_io_to_pes_2_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_36_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_36_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_36_io_to_pes_3_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_36_io_to_pes_3_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_36_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_36_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_36_io_to_pes_4_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_36_io_to_pes_4_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_36_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_36_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_36_io_to_pes_5_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_36_io_to_pes_5_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_36_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_36_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_36_io_to_pes_6_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_36_io_to_pes_6_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_36_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_36_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_36_io_to_pes_7_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_36_io_to_pes_7_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_36_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_36_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_36_io_to_pes_8_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_36_io_to_pes_8_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_36_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_36_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_36_io_to_pes_9_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_36_io_to_pes_9_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_36_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_36_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_36_io_to_pes_10_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_36_io_to_pes_10_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_36_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_36_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_36_io_to_pes_11_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_36_io_to_pes_11_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_36_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_36_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_36_io_to_pes_12_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_36_io_to_pes_12_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_36_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_36_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_36_io_to_pes_13_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_36_io_to_pes_13_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_36_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_36_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_36_io_to_pes_14_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_36_io_to_pes_14_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_36_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_36_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_36_io_to_pes_15_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_36_io_to_pes_15_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_36_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_36_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_36_io_to_pes_16_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_36_io_to_pes_16_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_36_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_36_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_36_io_to_pes_17_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_36_io_to_pes_17_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_36_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_36_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_36_io_to_pes_18_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_36_io_to_pes_18_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_36_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_36_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_36_io_to_pes_19_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_36_io_to_pes_19_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_36_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_36_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_36_io_to_pes_20_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_36_io_to_pes_20_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_36_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_36_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_36_io_to_pes_21_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_36_io_to_pes_21_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_36_io_to_mem_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_36_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_37_io_to_pes_0_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_37_io_to_pes_0_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_37_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_37_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_37_io_to_pes_1_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_37_io_to_pes_1_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_37_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_37_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_37_io_to_pes_2_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_37_io_to_pes_2_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_37_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_37_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_37_io_to_pes_3_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_37_io_to_pes_3_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_37_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_37_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_37_io_to_pes_4_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_37_io_to_pes_4_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_37_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_37_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_37_io_to_pes_5_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_37_io_to_pes_5_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_37_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_37_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_37_io_to_pes_6_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_37_io_to_pes_6_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_37_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_37_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_37_io_to_pes_7_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_37_io_to_pes_7_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_37_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_37_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_37_io_to_pes_8_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_37_io_to_pes_8_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_37_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_37_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_37_io_to_pes_9_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_37_io_to_pes_9_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_37_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_37_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_37_io_to_pes_10_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_37_io_to_pes_10_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_37_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_37_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_37_io_to_pes_11_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_37_io_to_pes_11_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_37_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_37_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_37_io_to_pes_12_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_37_io_to_pes_12_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_37_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_37_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_37_io_to_pes_13_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_37_io_to_pes_13_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_37_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_37_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_37_io_to_pes_14_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_37_io_to_pes_14_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_37_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_37_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_37_io_to_pes_15_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_37_io_to_pes_15_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_37_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_37_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_37_io_to_pes_16_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_37_io_to_pes_16_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_37_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_37_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_37_io_to_pes_17_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_37_io_to_pes_17_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_37_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_37_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_37_io_to_pes_18_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_37_io_to_pes_18_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_37_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_37_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_37_io_to_pes_19_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_37_io_to_pes_19_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_37_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_37_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_37_io_to_pes_20_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_37_io_to_pes_20_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_37_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_37_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_37_io_to_pes_21_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_37_io_to_pes_21_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_37_io_to_mem_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_37_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_38_io_to_pes_0_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_38_io_to_pes_0_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_38_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_38_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_38_io_to_pes_1_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_38_io_to_pes_1_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_38_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_38_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_38_io_to_pes_2_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_38_io_to_pes_2_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_38_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_38_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_38_io_to_pes_3_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_38_io_to_pes_3_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_38_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_38_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_38_io_to_pes_4_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_38_io_to_pes_4_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_38_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_38_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_38_io_to_pes_5_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_38_io_to_pes_5_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_38_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_38_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_38_io_to_pes_6_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_38_io_to_pes_6_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_38_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_38_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_38_io_to_pes_7_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_38_io_to_pes_7_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_38_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_38_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_38_io_to_pes_8_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_38_io_to_pes_8_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_38_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_38_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_38_io_to_pes_9_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_38_io_to_pes_9_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_38_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_38_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_38_io_to_pes_10_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_38_io_to_pes_10_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_38_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_38_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_38_io_to_pes_11_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_38_io_to_pes_11_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_38_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_38_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_38_io_to_pes_12_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_38_io_to_pes_12_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_38_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_38_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_38_io_to_pes_13_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_38_io_to_pes_13_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_38_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_38_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_38_io_to_pes_14_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_38_io_to_pes_14_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_38_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_38_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_38_io_to_pes_15_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_38_io_to_pes_15_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_38_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_38_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_38_io_to_pes_16_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_38_io_to_pes_16_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_38_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_38_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_38_io_to_pes_17_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_38_io_to_pes_17_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_38_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_38_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_38_io_to_pes_18_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_38_io_to_pes_18_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_38_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_38_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_38_io_to_pes_19_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_38_io_to_pes_19_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_38_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_38_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_38_io_to_pes_20_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_38_io_to_pes_20_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_38_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_38_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_38_io_to_pes_21_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_38_io_to_pes_21_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_38_io_to_mem_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_38_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_39_io_to_pes_0_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_39_io_to_pes_0_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_39_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_39_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_39_io_to_pes_1_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_39_io_to_pes_1_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_39_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_39_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_39_io_to_pes_2_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_39_io_to_pes_2_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_39_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_39_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_39_io_to_pes_3_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_39_io_to_pes_3_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_39_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_39_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_39_io_to_pes_4_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_39_io_to_pes_4_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_39_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_39_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_39_io_to_pes_5_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_39_io_to_pes_5_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_39_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_39_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_39_io_to_pes_6_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_39_io_to_pes_6_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_39_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_39_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_39_io_to_pes_7_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_39_io_to_pes_7_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_39_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_39_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_39_io_to_pes_8_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_39_io_to_pes_8_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_39_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_39_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_39_io_to_pes_9_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_39_io_to_pes_9_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_39_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_39_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_39_io_to_pes_10_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_39_io_to_pes_10_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_39_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_39_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_39_io_to_pes_11_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_39_io_to_pes_11_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_39_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_39_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_39_io_to_pes_12_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_39_io_to_pes_12_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_39_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_39_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_39_io_to_pes_13_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_39_io_to_pes_13_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_39_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_39_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_39_io_to_pes_14_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_39_io_to_pes_14_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_39_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_39_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_39_io_to_pes_15_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_39_io_to_pes_15_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_39_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_39_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_39_io_to_pes_16_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_39_io_to_pes_16_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_39_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_39_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_39_io_to_pes_17_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_39_io_to_pes_17_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_39_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_39_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_39_io_to_pes_18_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_39_io_to_pes_18_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_39_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_39_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_39_io_to_pes_19_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_39_io_to_pes_19_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_39_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_39_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_39_io_to_pes_20_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_39_io_to_pes_20_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_39_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_39_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_39_io_to_pes_21_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_39_io_to_pes_21_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_39_io_to_mem_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_39_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_40_io_to_pes_0_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_40_io_to_pes_0_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_40_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_40_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_40_io_to_pes_1_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_40_io_to_pes_1_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_40_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_40_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_40_io_to_pes_2_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_40_io_to_pes_2_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_40_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_40_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_40_io_to_pes_3_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_40_io_to_pes_3_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_40_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_40_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_40_io_to_pes_4_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_40_io_to_pes_4_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_40_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_40_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_40_io_to_pes_5_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_40_io_to_pes_5_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_40_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_40_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_40_io_to_pes_6_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_40_io_to_pes_6_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_40_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_40_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_40_io_to_pes_7_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_40_io_to_pes_7_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_40_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_40_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_40_io_to_pes_8_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_40_io_to_pes_8_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_40_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_40_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_40_io_to_pes_9_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_40_io_to_pes_9_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_40_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_40_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_40_io_to_pes_10_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_40_io_to_pes_10_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_40_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_40_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_40_io_to_pes_11_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_40_io_to_pes_11_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_40_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_40_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_40_io_to_pes_12_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_40_io_to_pes_12_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_40_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_40_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_40_io_to_pes_13_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_40_io_to_pes_13_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_40_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_40_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_40_io_to_pes_14_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_40_io_to_pes_14_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_40_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_40_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_40_io_to_pes_15_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_40_io_to_pes_15_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_40_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_40_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_40_io_to_pes_16_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_40_io_to_pes_16_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_40_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_40_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_40_io_to_pes_17_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_40_io_to_pes_17_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_40_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_40_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_40_io_to_pes_18_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_40_io_to_pes_18_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_40_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_40_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_40_io_to_pes_19_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_40_io_to_pes_19_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_40_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_40_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_40_io_to_pes_20_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_40_io_to_pes_20_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_40_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_40_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_40_io_to_pes_21_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_40_io_to_pes_21_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_40_io_to_mem_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_40_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_41_io_to_pes_0_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_41_io_to_pes_0_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_41_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_41_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_41_io_to_pes_1_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_41_io_to_pes_1_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_41_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_41_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_41_io_to_pes_2_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_41_io_to_pes_2_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_41_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_41_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_41_io_to_pes_3_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_41_io_to_pes_3_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_41_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_41_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_41_io_to_pes_4_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_41_io_to_pes_4_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_41_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_41_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_41_io_to_pes_5_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_41_io_to_pes_5_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_41_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_41_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_41_io_to_pes_6_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_41_io_to_pes_6_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_41_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_41_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_41_io_to_pes_7_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_41_io_to_pes_7_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_41_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_41_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_41_io_to_pes_8_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_41_io_to_pes_8_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_41_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_41_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_41_io_to_pes_9_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_41_io_to_pes_9_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_41_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_41_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_41_io_to_pes_10_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_41_io_to_pes_10_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_41_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_41_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_41_io_to_pes_11_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_41_io_to_pes_11_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_41_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_41_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_41_io_to_pes_12_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_41_io_to_pes_12_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_41_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_41_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_41_io_to_pes_13_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_41_io_to_pes_13_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_41_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_41_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_41_io_to_pes_14_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_41_io_to_pes_14_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_41_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_41_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_41_io_to_pes_15_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_41_io_to_pes_15_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_41_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_41_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_41_io_to_pes_16_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_41_io_to_pes_16_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_41_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_41_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_41_io_to_pes_17_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_41_io_to_pes_17_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_41_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_41_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_41_io_to_pes_18_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_41_io_to_pes_18_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_41_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_41_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_41_io_to_pes_19_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_41_io_to_pes_19_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_41_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_41_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_41_io_to_pes_20_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_41_io_to_pes_20_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_41_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_41_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_41_io_to_pes_21_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_41_io_to_pes_21_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_41_io_to_mem_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_41_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_42_io_to_pes_0_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_42_io_to_pes_0_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_42_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_42_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_42_io_to_pes_1_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_42_io_to_pes_1_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_42_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_42_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_42_io_to_pes_2_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_42_io_to_pes_2_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_42_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_42_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_42_io_to_pes_3_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_42_io_to_pes_3_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_42_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_42_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_42_io_to_pes_4_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_42_io_to_pes_4_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_42_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_42_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_42_io_to_pes_5_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_42_io_to_pes_5_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_42_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_42_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_42_io_to_pes_6_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_42_io_to_pes_6_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_42_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_42_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_42_io_to_pes_7_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_42_io_to_pes_7_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_42_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_42_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_42_io_to_pes_8_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_42_io_to_pes_8_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_42_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_42_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_42_io_to_pes_9_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_42_io_to_pes_9_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_42_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_42_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_42_io_to_pes_10_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_42_io_to_pes_10_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_42_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_42_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_42_io_to_pes_11_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_42_io_to_pes_11_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_42_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_42_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_42_io_to_pes_12_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_42_io_to_pes_12_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_42_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_42_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_42_io_to_pes_13_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_42_io_to_pes_13_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_42_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_42_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_42_io_to_pes_14_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_42_io_to_pes_14_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_42_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_42_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_42_io_to_pes_15_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_42_io_to_pes_15_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_42_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_42_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_42_io_to_pes_16_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_42_io_to_pes_16_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_42_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_42_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_42_io_to_pes_17_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_42_io_to_pes_17_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_42_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_42_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_42_io_to_pes_18_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_42_io_to_pes_18_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_42_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_42_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_42_io_to_pes_19_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_42_io_to_pes_19_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_42_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_42_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_42_io_to_pes_20_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_42_io_to_pes_20_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_42_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_42_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_42_io_to_pes_21_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_42_io_to_pes_21_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_42_io_to_mem_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_42_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_43_io_to_pes_0_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_43_io_to_pes_0_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_43_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_43_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_43_io_to_pes_1_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_43_io_to_pes_1_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_43_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_43_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_43_io_to_pes_2_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_43_io_to_pes_2_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_43_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_43_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_43_io_to_pes_3_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_43_io_to_pes_3_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_43_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_43_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_43_io_to_pes_4_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_43_io_to_pes_4_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_43_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_43_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_43_io_to_pes_5_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_43_io_to_pes_5_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_43_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_43_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_43_io_to_pes_6_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_43_io_to_pes_6_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_43_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_43_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_43_io_to_pes_7_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_43_io_to_pes_7_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_43_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_43_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_43_io_to_pes_8_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_43_io_to_pes_8_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_43_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_43_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_43_io_to_pes_9_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_43_io_to_pes_9_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_43_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_43_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_43_io_to_pes_10_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_43_io_to_pes_10_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_43_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_43_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_43_io_to_pes_11_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_43_io_to_pes_11_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_43_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_43_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_43_io_to_pes_12_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_43_io_to_pes_12_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_43_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_43_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_43_io_to_pes_13_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_43_io_to_pes_13_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_43_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_43_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_43_io_to_pes_14_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_43_io_to_pes_14_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_43_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_43_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_43_io_to_pes_15_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_43_io_to_pes_15_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_43_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_43_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_43_io_to_pes_16_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_43_io_to_pes_16_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_43_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_43_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_43_io_to_pes_17_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_43_io_to_pes_17_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_43_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_43_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_43_io_to_pes_18_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_43_io_to_pes_18_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_43_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_43_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_43_io_to_pes_19_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_43_io_to_pes_19_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_43_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_43_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_43_io_to_pes_20_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_43_io_to_pes_20_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_43_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_43_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_43_io_to_pes_21_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_43_io_to_pes_21_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_43_io_to_mem_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_43_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_44_io_to_pes_0_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_44_io_to_pes_0_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_44_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_44_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_44_io_to_pes_1_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_44_io_to_pes_1_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_44_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_44_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_44_io_to_pes_2_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_44_io_to_pes_2_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_44_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_44_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_44_io_to_pes_3_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_44_io_to_pes_3_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_44_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_44_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_44_io_to_pes_4_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_44_io_to_pes_4_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_44_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_44_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_44_io_to_pes_5_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_44_io_to_pes_5_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_44_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_44_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_44_io_to_pes_6_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_44_io_to_pes_6_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_44_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_44_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_44_io_to_pes_7_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_44_io_to_pes_7_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_44_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_44_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_44_io_to_pes_8_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_44_io_to_pes_8_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_44_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_44_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_44_io_to_pes_9_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_44_io_to_pes_9_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_44_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_44_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_44_io_to_pes_10_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_44_io_to_pes_10_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_44_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_44_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_44_io_to_pes_11_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_44_io_to_pes_11_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_44_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_44_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_44_io_to_pes_12_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_44_io_to_pes_12_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_44_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_44_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_44_io_to_pes_13_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_44_io_to_pes_13_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_44_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_44_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_44_io_to_pes_14_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_44_io_to_pes_14_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_44_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_44_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_44_io_to_pes_15_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_44_io_to_pes_15_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_44_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_44_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_44_io_to_pes_16_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_44_io_to_pes_16_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_44_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_44_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_44_io_to_pes_17_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_44_io_to_pes_17_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_44_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_44_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_44_io_to_pes_18_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_44_io_to_pes_18_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_44_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_44_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_44_io_to_pes_19_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_44_io_to_pes_19_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_44_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_44_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_44_io_to_pes_20_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_44_io_to_pes_20_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_44_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_44_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_44_io_to_pes_21_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_44_io_to_pes_21_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_44_io_to_mem_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_44_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_45_io_to_pes_0_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_45_io_to_pes_0_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_45_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_45_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_45_io_to_pes_1_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_45_io_to_pes_1_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_45_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_45_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_45_io_to_pes_2_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_45_io_to_pes_2_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_45_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_45_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_45_io_to_pes_3_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_45_io_to_pes_3_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_45_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_45_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_45_io_to_pes_4_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_45_io_to_pes_4_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_45_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_45_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_45_io_to_pes_5_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_45_io_to_pes_5_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_45_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_45_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_45_io_to_pes_6_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_45_io_to_pes_6_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_45_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_45_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_45_io_to_pes_7_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_45_io_to_pes_7_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_45_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_45_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_45_io_to_pes_8_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_45_io_to_pes_8_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_45_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_45_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_45_io_to_pes_9_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_45_io_to_pes_9_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_45_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_45_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_45_io_to_pes_10_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_45_io_to_pes_10_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_45_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_45_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_45_io_to_pes_11_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_45_io_to_pes_11_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_45_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_45_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_45_io_to_pes_12_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_45_io_to_pes_12_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_45_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_45_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_45_io_to_pes_13_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_45_io_to_pes_13_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_45_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_45_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_45_io_to_pes_14_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_45_io_to_pes_14_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_45_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_45_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_45_io_to_pes_15_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_45_io_to_pes_15_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_45_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_45_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_45_io_to_pes_16_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_45_io_to_pes_16_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_45_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_45_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_45_io_to_pes_17_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_45_io_to_pes_17_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_45_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_45_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_45_io_to_pes_18_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_45_io_to_pes_18_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_45_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_45_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_45_io_to_pes_19_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_45_io_to_pes_19_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_45_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_45_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_45_io_to_pes_20_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_45_io_to_pes_20_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_45_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_45_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_45_io_to_pes_21_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_45_io_to_pes_21_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_45_io_to_mem_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_45_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_46_io_to_pes_0_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_46_io_to_pes_0_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_46_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_46_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_46_io_to_pes_1_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_46_io_to_pes_1_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_46_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_46_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_46_io_to_pes_2_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_46_io_to_pes_2_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_46_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_46_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_46_io_to_pes_3_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_46_io_to_pes_3_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_46_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_46_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_46_io_to_pes_4_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_46_io_to_pes_4_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_46_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_46_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_46_io_to_pes_5_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_46_io_to_pes_5_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_46_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_46_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_46_io_to_pes_6_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_46_io_to_pes_6_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_46_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_46_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_46_io_to_pes_7_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_46_io_to_pes_7_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_46_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_46_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_46_io_to_pes_8_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_46_io_to_pes_8_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_46_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_46_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_46_io_to_pes_9_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_46_io_to_pes_9_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_46_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_46_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_46_io_to_pes_10_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_46_io_to_pes_10_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_46_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_46_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_46_io_to_pes_11_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_46_io_to_pes_11_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_46_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_46_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_46_io_to_pes_12_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_46_io_to_pes_12_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_46_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_46_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_46_io_to_pes_13_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_46_io_to_pes_13_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_46_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_46_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_46_io_to_pes_14_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_46_io_to_pes_14_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_46_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_46_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_46_io_to_pes_15_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_46_io_to_pes_15_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_46_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_46_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_46_io_to_pes_16_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_46_io_to_pes_16_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_46_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_46_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_46_io_to_pes_17_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_46_io_to_pes_17_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_46_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_46_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_46_io_to_pes_18_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_46_io_to_pes_18_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_46_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_46_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_46_io_to_pes_19_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_46_io_to_pes_19_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_46_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_46_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_46_io_to_pes_20_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_46_io_to_pes_20_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_46_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_46_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_46_io_to_pes_21_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_46_io_to_pes_21_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_46_io_to_mem_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_46_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_47_io_to_pes_0_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_47_io_to_pes_0_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_47_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_47_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_47_io_to_pes_1_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_47_io_to_pes_1_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_47_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_47_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_47_io_to_pes_2_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_47_io_to_pes_2_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_47_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_47_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_47_io_to_pes_3_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_47_io_to_pes_3_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_47_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_47_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_47_io_to_pes_4_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_47_io_to_pes_4_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_47_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_47_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_47_io_to_pes_5_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_47_io_to_pes_5_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_47_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_47_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_47_io_to_pes_6_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_47_io_to_pes_6_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_47_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_47_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_47_io_to_pes_7_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_47_io_to_pes_7_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_47_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_47_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_47_io_to_pes_8_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_47_io_to_pes_8_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_47_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_47_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_47_io_to_pes_9_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_47_io_to_pes_9_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_47_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_47_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_47_io_to_pes_10_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_47_io_to_pes_10_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_47_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_47_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_47_io_to_pes_11_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_47_io_to_pes_11_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_47_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_47_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_47_io_to_pes_12_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_47_io_to_pes_12_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_47_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_47_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_47_io_to_pes_13_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_47_io_to_pes_13_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_47_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_47_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_47_io_to_pes_14_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_47_io_to_pes_14_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_47_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_47_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_47_io_to_pes_15_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_47_io_to_pes_15_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_47_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_47_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_47_io_to_pes_16_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_47_io_to_pes_16_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_47_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_47_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_47_io_to_pes_17_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_47_io_to_pes_17_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_47_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_47_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_47_io_to_pes_18_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_47_io_to_pes_18_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_47_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_47_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_47_io_to_pes_19_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_47_io_to_pes_19_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_47_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_47_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_47_io_to_pes_20_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_47_io_to_pes_20_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_47_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_47_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_47_io_to_pes_21_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_47_io_to_pes_21_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_47_io_to_mem_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_47_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_48_io_to_pes_0_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_48_io_to_pes_0_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_48_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_48_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_48_io_to_pes_1_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_48_io_to_pes_1_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_48_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_48_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_48_io_to_pes_2_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_48_io_to_pes_2_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_48_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_48_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_48_io_to_pes_3_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_48_io_to_pes_3_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_48_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_48_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_48_io_to_pes_4_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_48_io_to_pes_4_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_48_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_48_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_48_io_to_pes_5_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_48_io_to_pes_5_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_48_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_48_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_48_io_to_pes_6_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_48_io_to_pes_6_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_48_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_48_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_48_io_to_pes_7_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_48_io_to_pes_7_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_48_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_48_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_48_io_to_pes_8_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_48_io_to_pes_8_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_48_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_48_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_48_io_to_pes_9_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_48_io_to_pes_9_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_48_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_48_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_48_io_to_pes_10_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_48_io_to_pes_10_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_48_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_48_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_48_io_to_pes_11_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_48_io_to_pes_11_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_48_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_48_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_48_io_to_pes_12_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_48_io_to_pes_12_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_48_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_48_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_48_io_to_pes_13_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_48_io_to_pes_13_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_48_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_48_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_48_io_to_pes_14_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_48_io_to_pes_14_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_48_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_48_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_48_io_to_pes_15_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_48_io_to_pes_15_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_48_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_48_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_48_io_to_pes_16_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_48_io_to_pes_16_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_48_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_48_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_48_io_to_pes_17_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_48_io_to_pes_17_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_48_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_48_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_48_io_to_pes_18_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_48_io_to_pes_18_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_48_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_48_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_48_io_to_pes_19_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_48_io_to_pes_19_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_48_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_48_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_48_io_to_pes_20_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_48_io_to_pes_20_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_48_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_48_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_48_io_to_pes_21_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_48_io_to_pes_21_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_48_io_to_mem_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_48_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_49_io_to_pes_0_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_49_io_to_pes_0_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_49_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_49_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_49_io_to_pes_1_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_49_io_to_pes_1_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_49_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_49_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_49_io_to_pes_2_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_49_io_to_pes_2_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_49_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_49_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_49_io_to_pes_3_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_49_io_to_pes_3_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_49_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_49_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_49_io_to_pes_4_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_49_io_to_pes_4_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_49_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_49_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_49_io_to_pes_5_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_49_io_to_pes_5_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_49_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_49_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_49_io_to_pes_6_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_49_io_to_pes_6_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_49_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_49_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_49_io_to_pes_7_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_49_io_to_pes_7_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_49_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_49_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_49_io_to_pes_8_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_49_io_to_pes_8_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_49_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_49_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_49_io_to_pes_9_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_49_io_to_pes_9_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_49_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_49_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_49_io_to_pes_10_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_49_io_to_pes_10_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_49_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_49_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_49_io_to_pes_11_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_49_io_to_pes_11_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_49_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_49_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_49_io_to_pes_12_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_49_io_to_pes_12_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_49_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_49_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_49_io_to_pes_13_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_49_io_to_pes_13_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_49_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_49_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_49_io_to_pes_14_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_49_io_to_pes_14_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_49_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_49_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_49_io_to_pes_15_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_49_io_to_pes_15_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_49_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_49_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_49_io_to_pes_16_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_49_io_to_pes_16_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_49_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_49_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_49_io_to_pes_17_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_49_io_to_pes_17_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_49_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_49_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_49_io_to_pes_18_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_49_io_to_pes_18_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_49_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_49_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_49_io_to_pes_19_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_49_io_to_pes_19_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_49_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_49_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_49_io_to_pes_20_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_49_io_to_pes_20_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_49_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_49_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_49_io_to_pes_21_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_49_io_to_pes_21_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_49_io_to_mem_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_49_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_50_io_to_pes_0_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_50_io_to_pes_0_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_50_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_50_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_50_io_to_pes_1_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_50_io_to_pes_1_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_50_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_50_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_50_io_to_pes_2_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_50_io_to_pes_2_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_50_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_50_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_50_io_to_pes_3_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_50_io_to_pes_3_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_50_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_50_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_50_io_to_pes_4_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_50_io_to_pes_4_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_50_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_50_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_50_io_to_pes_5_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_50_io_to_pes_5_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_50_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_50_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_50_io_to_pes_6_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_50_io_to_pes_6_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_50_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_50_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_50_io_to_pes_7_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_50_io_to_pes_7_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_50_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_50_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_50_io_to_pes_8_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_50_io_to_pes_8_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_50_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_50_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_50_io_to_pes_9_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_50_io_to_pes_9_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_50_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_50_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_50_io_to_pes_10_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_50_io_to_pes_10_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_50_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_50_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_50_io_to_pes_11_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_50_io_to_pes_11_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_50_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_50_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_50_io_to_pes_12_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_50_io_to_pes_12_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_50_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_50_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_50_io_to_pes_13_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_50_io_to_pes_13_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_50_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_50_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_50_io_to_pes_14_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_50_io_to_pes_14_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_50_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_50_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_50_io_to_pes_15_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_50_io_to_pes_15_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_50_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_50_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_50_io_to_pes_16_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_50_io_to_pes_16_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_50_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_50_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_50_io_to_pes_17_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_50_io_to_pes_17_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_50_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_50_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_50_io_to_pes_18_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_50_io_to_pes_18_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_50_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_50_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_50_io_to_pes_19_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_50_io_to_pes_19_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_50_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_50_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_50_io_to_pes_20_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_50_io_to_pes_20_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_50_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_50_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_50_io_to_pes_21_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_50_io_to_pes_21_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_50_io_to_mem_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_50_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_51_io_to_pes_0_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_51_io_to_pes_0_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_51_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_51_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_51_io_to_pes_1_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_51_io_to_pes_1_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_51_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_51_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_51_io_to_pes_2_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_51_io_to_pes_2_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_51_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_51_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_51_io_to_pes_3_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_51_io_to_pes_3_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_51_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_51_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_51_io_to_pes_4_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_51_io_to_pes_4_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_51_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_51_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_51_io_to_pes_5_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_51_io_to_pes_5_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_51_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_51_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_51_io_to_pes_6_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_51_io_to_pes_6_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_51_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_51_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_51_io_to_pes_7_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_51_io_to_pes_7_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_51_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_51_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_51_io_to_pes_8_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_51_io_to_pes_8_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_51_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_51_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_51_io_to_pes_9_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_51_io_to_pes_9_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_51_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_51_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_51_io_to_pes_10_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_51_io_to_pes_10_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_51_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_51_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_51_io_to_pes_11_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_51_io_to_pes_11_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_51_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_51_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_51_io_to_pes_12_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_51_io_to_pes_12_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_51_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_51_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_51_io_to_pes_13_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_51_io_to_pes_13_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_51_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_51_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_51_io_to_pes_14_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_51_io_to_pes_14_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_51_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_51_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_51_io_to_pes_15_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_51_io_to_pes_15_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_51_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_51_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_51_io_to_pes_16_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_51_io_to_pes_16_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_51_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_51_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_51_io_to_pes_17_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_51_io_to_pes_17_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_51_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_51_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_51_io_to_pes_18_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_51_io_to_pes_18_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_51_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_51_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_51_io_to_pes_19_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_51_io_to_pes_19_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_51_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_51_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_51_io_to_pes_20_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_51_io_to_pes_20_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_51_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_51_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_51_io_to_pes_21_in_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_51_io_to_pes_21_in_bits; // @[pe.scala 229:13]
  wire  PENetwork_51_io_to_mem_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_51_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_52_clock; // @[pe.scala 229:13]
  wire  PENetwork_52_reset; // @[pe.scala 229:13]
  wire  PENetwork_52_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_52_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_52_io_to_pes_0_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_52_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_52_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_52_io_to_pes_1_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_52_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_52_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_52_io_to_pes_2_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_52_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_52_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_52_io_to_pes_3_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_52_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_52_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_52_io_to_pes_4_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_52_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_52_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_52_io_to_pes_5_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_52_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_52_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_52_io_to_pes_6_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_52_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_52_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_52_io_to_pes_7_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_52_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_52_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_52_io_to_pes_8_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_52_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_52_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_52_io_to_pes_9_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_52_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_52_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_52_io_to_pes_10_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_52_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_52_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_52_io_to_pes_11_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_52_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_52_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_52_io_to_pes_12_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_52_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_52_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_52_io_to_pes_13_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_52_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_52_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_52_io_to_pes_14_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_52_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_52_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_52_io_to_pes_15_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_52_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_52_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_52_io_to_pes_16_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_52_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_52_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_52_io_to_pes_17_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_52_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_52_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_52_io_to_pes_18_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_52_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_52_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_52_io_to_pes_19_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_52_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_52_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_52_io_to_pes_20_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_52_io_to_pes_21_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_52_io_to_pes_21_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_52_io_to_pes_21_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_52_io_to_mem_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_52_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_52_io_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_53_clock; // @[pe.scala 229:13]
  wire  PENetwork_53_reset; // @[pe.scala 229:13]
  wire  PENetwork_53_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_53_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_53_io_to_pes_0_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_53_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_53_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_53_io_to_pes_1_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_53_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_53_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_53_io_to_pes_2_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_53_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_53_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_53_io_to_pes_3_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_53_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_53_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_53_io_to_pes_4_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_53_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_53_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_53_io_to_pes_5_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_53_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_53_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_53_io_to_pes_6_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_53_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_53_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_53_io_to_pes_7_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_53_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_53_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_53_io_to_pes_8_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_53_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_53_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_53_io_to_pes_9_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_53_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_53_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_53_io_to_pes_10_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_53_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_53_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_53_io_to_pes_11_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_53_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_53_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_53_io_to_pes_12_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_53_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_53_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_53_io_to_pes_13_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_53_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_53_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_53_io_to_pes_14_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_53_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_53_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_53_io_to_pes_15_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_53_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_53_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_53_io_to_pes_16_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_53_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_53_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_53_io_to_pes_17_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_53_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_53_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_53_io_to_pes_18_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_53_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_53_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_53_io_to_pes_19_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_53_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_53_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_53_io_to_pes_20_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_53_io_to_pes_21_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_53_io_to_pes_21_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_53_io_to_pes_21_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_53_io_to_mem_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_53_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_53_io_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_54_clock; // @[pe.scala 229:13]
  wire  PENetwork_54_reset; // @[pe.scala 229:13]
  wire  PENetwork_54_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_54_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_54_io_to_pes_0_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_54_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_54_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_54_io_to_pes_1_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_54_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_54_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_54_io_to_pes_2_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_54_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_54_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_54_io_to_pes_3_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_54_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_54_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_54_io_to_pes_4_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_54_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_54_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_54_io_to_pes_5_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_54_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_54_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_54_io_to_pes_6_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_54_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_54_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_54_io_to_pes_7_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_54_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_54_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_54_io_to_pes_8_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_54_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_54_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_54_io_to_pes_9_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_54_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_54_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_54_io_to_pes_10_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_54_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_54_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_54_io_to_pes_11_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_54_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_54_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_54_io_to_pes_12_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_54_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_54_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_54_io_to_pes_13_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_54_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_54_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_54_io_to_pes_14_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_54_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_54_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_54_io_to_pes_15_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_54_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_54_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_54_io_to_pes_16_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_54_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_54_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_54_io_to_pes_17_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_54_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_54_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_54_io_to_pes_18_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_54_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_54_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_54_io_to_pes_19_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_54_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_54_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_54_io_to_pes_20_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_54_io_to_pes_21_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_54_io_to_pes_21_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_54_io_to_pes_21_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_54_io_to_mem_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_54_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_54_io_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_55_clock; // @[pe.scala 229:13]
  wire  PENetwork_55_reset; // @[pe.scala 229:13]
  wire  PENetwork_55_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_55_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_55_io_to_pes_0_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_55_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_55_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_55_io_to_pes_1_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_55_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_55_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_55_io_to_pes_2_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_55_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_55_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_55_io_to_pes_3_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_55_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_55_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_55_io_to_pes_4_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_55_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_55_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_55_io_to_pes_5_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_55_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_55_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_55_io_to_pes_6_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_55_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_55_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_55_io_to_pes_7_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_55_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_55_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_55_io_to_pes_8_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_55_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_55_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_55_io_to_pes_9_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_55_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_55_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_55_io_to_pes_10_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_55_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_55_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_55_io_to_pes_11_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_55_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_55_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_55_io_to_pes_12_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_55_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_55_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_55_io_to_pes_13_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_55_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_55_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_55_io_to_pes_14_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_55_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_55_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_55_io_to_pes_15_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_55_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_55_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_55_io_to_pes_16_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_55_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_55_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_55_io_to_pes_17_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_55_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_55_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_55_io_to_pes_18_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_55_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_55_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_55_io_to_pes_19_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_55_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_55_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_55_io_to_pes_20_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_55_io_to_pes_21_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_55_io_to_pes_21_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_55_io_to_pes_21_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_55_io_to_mem_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_55_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_55_io_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_56_clock; // @[pe.scala 229:13]
  wire  PENetwork_56_reset; // @[pe.scala 229:13]
  wire  PENetwork_56_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_56_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_56_io_to_pes_0_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_56_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_56_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_56_io_to_pes_1_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_56_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_56_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_56_io_to_pes_2_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_56_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_56_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_56_io_to_pes_3_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_56_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_56_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_56_io_to_pes_4_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_56_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_56_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_56_io_to_pes_5_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_56_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_56_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_56_io_to_pes_6_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_56_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_56_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_56_io_to_pes_7_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_56_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_56_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_56_io_to_pes_8_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_56_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_56_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_56_io_to_pes_9_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_56_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_56_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_56_io_to_pes_10_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_56_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_56_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_56_io_to_pes_11_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_56_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_56_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_56_io_to_pes_12_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_56_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_56_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_56_io_to_pes_13_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_56_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_56_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_56_io_to_pes_14_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_56_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_56_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_56_io_to_pes_15_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_56_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_56_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_56_io_to_pes_16_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_56_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_56_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_56_io_to_pes_17_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_56_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_56_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_56_io_to_pes_18_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_56_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_56_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_56_io_to_pes_19_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_56_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_56_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_56_io_to_pes_20_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_56_io_to_pes_21_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_56_io_to_pes_21_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_56_io_to_pes_21_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_56_io_to_mem_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_56_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_56_io_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_57_clock; // @[pe.scala 229:13]
  wire  PENetwork_57_reset; // @[pe.scala 229:13]
  wire  PENetwork_57_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_57_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_57_io_to_pes_0_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_57_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_57_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_57_io_to_pes_1_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_57_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_57_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_57_io_to_pes_2_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_57_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_57_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_57_io_to_pes_3_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_57_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_57_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_57_io_to_pes_4_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_57_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_57_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_57_io_to_pes_5_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_57_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_57_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_57_io_to_pes_6_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_57_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_57_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_57_io_to_pes_7_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_57_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_57_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_57_io_to_pes_8_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_57_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_57_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_57_io_to_pes_9_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_57_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_57_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_57_io_to_pes_10_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_57_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_57_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_57_io_to_pes_11_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_57_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_57_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_57_io_to_pes_12_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_57_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_57_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_57_io_to_pes_13_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_57_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_57_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_57_io_to_pes_14_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_57_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_57_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_57_io_to_pes_15_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_57_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_57_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_57_io_to_pes_16_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_57_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_57_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_57_io_to_pes_17_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_57_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_57_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_57_io_to_pes_18_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_57_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_57_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_57_io_to_pes_19_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_57_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_57_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_57_io_to_pes_20_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_57_io_to_pes_21_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_57_io_to_pes_21_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_57_io_to_pes_21_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_57_io_to_mem_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_57_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_57_io_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_58_clock; // @[pe.scala 229:13]
  wire  PENetwork_58_reset; // @[pe.scala 229:13]
  wire  PENetwork_58_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_58_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_58_io_to_pes_0_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_58_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_58_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_58_io_to_pes_1_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_58_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_58_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_58_io_to_pes_2_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_58_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_58_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_58_io_to_pes_3_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_58_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_58_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_58_io_to_pes_4_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_58_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_58_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_58_io_to_pes_5_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_58_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_58_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_58_io_to_pes_6_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_58_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_58_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_58_io_to_pes_7_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_58_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_58_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_58_io_to_pes_8_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_58_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_58_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_58_io_to_pes_9_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_58_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_58_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_58_io_to_pes_10_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_58_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_58_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_58_io_to_pes_11_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_58_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_58_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_58_io_to_pes_12_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_58_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_58_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_58_io_to_pes_13_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_58_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_58_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_58_io_to_pes_14_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_58_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_58_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_58_io_to_pes_15_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_58_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_58_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_58_io_to_pes_16_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_58_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_58_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_58_io_to_pes_17_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_58_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_58_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_58_io_to_pes_18_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_58_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_58_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_58_io_to_pes_19_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_58_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_58_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_58_io_to_pes_20_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_58_io_to_pes_21_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_58_io_to_pes_21_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_58_io_to_pes_21_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_58_io_to_mem_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_58_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_58_io_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_59_clock; // @[pe.scala 229:13]
  wire  PENetwork_59_reset; // @[pe.scala 229:13]
  wire  PENetwork_59_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_59_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_59_io_to_pes_0_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_59_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_59_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_59_io_to_pes_1_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_59_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_59_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_59_io_to_pes_2_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_59_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_59_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_59_io_to_pes_3_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_59_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_59_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_59_io_to_pes_4_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_59_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_59_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_59_io_to_pes_5_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_59_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_59_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_59_io_to_pes_6_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_59_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_59_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_59_io_to_pes_7_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_59_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_59_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_59_io_to_pes_8_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_59_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_59_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_59_io_to_pes_9_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_59_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_59_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_59_io_to_pes_10_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_59_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_59_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_59_io_to_pes_11_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_59_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_59_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_59_io_to_pes_12_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_59_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_59_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_59_io_to_pes_13_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_59_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_59_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_59_io_to_pes_14_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_59_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_59_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_59_io_to_pes_15_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_59_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_59_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_59_io_to_pes_16_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_59_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_59_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_59_io_to_pes_17_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_59_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_59_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_59_io_to_pes_18_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_59_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_59_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_59_io_to_pes_19_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_59_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_59_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_59_io_to_pes_20_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_59_io_to_pes_21_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_59_io_to_pes_21_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_59_io_to_pes_21_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_59_io_to_mem_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_59_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_59_io_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_60_clock; // @[pe.scala 229:13]
  wire  PENetwork_60_reset; // @[pe.scala 229:13]
  wire  PENetwork_60_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_60_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_60_io_to_pes_0_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_60_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_60_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_60_io_to_pes_1_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_60_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_60_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_60_io_to_pes_2_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_60_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_60_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_60_io_to_pes_3_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_60_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_60_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_60_io_to_pes_4_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_60_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_60_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_60_io_to_pes_5_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_60_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_60_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_60_io_to_pes_6_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_60_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_60_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_60_io_to_pes_7_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_60_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_60_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_60_io_to_pes_8_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_60_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_60_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_60_io_to_pes_9_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_60_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_60_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_60_io_to_pes_10_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_60_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_60_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_60_io_to_pes_11_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_60_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_60_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_60_io_to_pes_12_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_60_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_60_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_60_io_to_pes_13_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_60_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_60_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_60_io_to_pes_14_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_60_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_60_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_60_io_to_pes_15_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_60_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_60_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_60_io_to_pes_16_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_60_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_60_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_60_io_to_pes_17_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_60_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_60_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_60_io_to_pes_18_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_60_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_60_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_60_io_to_pes_19_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_60_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_60_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_60_io_to_pes_20_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_60_io_to_pes_21_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_60_io_to_pes_21_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_60_io_to_pes_21_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_60_io_to_mem_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_60_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_60_io_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_61_clock; // @[pe.scala 229:13]
  wire  PENetwork_61_reset; // @[pe.scala 229:13]
  wire  PENetwork_61_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_61_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_61_io_to_pes_0_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_61_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_61_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_61_io_to_pes_1_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_61_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_61_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_61_io_to_pes_2_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_61_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_61_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_61_io_to_pes_3_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_61_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_61_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_61_io_to_pes_4_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_61_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_61_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_61_io_to_pes_5_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_61_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_61_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_61_io_to_pes_6_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_61_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_61_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_61_io_to_pes_7_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_61_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_61_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_61_io_to_pes_8_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_61_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_61_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_61_io_to_pes_9_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_61_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_61_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_61_io_to_pes_10_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_61_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_61_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_61_io_to_pes_11_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_61_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_61_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_61_io_to_pes_12_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_61_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_61_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_61_io_to_pes_13_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_61_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_61_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_61_io_to_pes_14_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_61_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_61_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_61_io_to_pes_15_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_61_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_61_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_61_io_to_pes_16_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_61_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_61_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_61_io_to_pes_17_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_61_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_61_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_61_io_to_pes_18_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_61_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_61_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_61_io_to_pes_19_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_61_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_61_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_61_io_to_pes_20_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_61_io_to_pes_21_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_61_io_to_pes_21_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_61_io_to_pes_21_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_61_io_to_mem_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_61_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_61_io_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_62_clock; // @[pe.scala 229:13]
  wire  PENetwork_62_reset; // @[pe.scala 229:13]
  wire  PENetwork_62_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_62_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_62_io_to_pes_0_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_62_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_62_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_62_io_to_pes_1_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_62_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_62_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_62_io_to_pes_2_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_62_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_62_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_62_io_to_pes_3_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_62_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_62_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_62_io_to_pes_4_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_62_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_62_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_62_io_to_pes_5_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_62_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_62_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_62_io_to_pes_6_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_62_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_62_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_62_io_to_pes_7_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_62_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_62_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_62_io_to_pes_8_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_62_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_62_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_62_io_to_pes_9_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_62_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_62_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_62_io_to_pes_10_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_62_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_62_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_62_io_to_pes_11_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_62_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_62_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_62_io_to_pes_12_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_62_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_62_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_62_io_to_pes_13_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_62_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_62_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_62_io_to_pes_14_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_62_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_62_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_62_io_to_pes_15_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_62_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_62_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_62_io_to_pes_16_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_62_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_62_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_62_io_to_pes_17_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_62_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_62_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_62_io_to_pes_18_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_62_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_62_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_62_io_to_pes_19_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_62_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_62_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_62_io_to_pes_20_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_62_io_to_pes_21_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_62_io_to_pes_21_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_62_io_to_pes_21_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_62_io_to_mem_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_62_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_62_io_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_63_clock; // @[pe.scala 229:13]
  wire  PENetwork_63_reset; // @[pe.scala 229:13]
  wire  PENetwork_63_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_63_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_63_io_to_pes_0_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_63_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_63_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_63_io_to_pes_1_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_63_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_63_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_63_io_to_pes_2_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_63_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_63_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_63_io_to_pes_3_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_63_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_63_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_63_io_to_pes_4_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_63_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_63_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_63_io_to_pes_5_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_63_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_63_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_63_io_to_pes_6_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_63_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_63_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_63_io_to_pes_7_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_63_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_63_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_63_io_to_pes_8_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_63_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_63_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_63_io_to_pes_9_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_63_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_63_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_63_io_to_pes_10_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_63_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_63_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_63_io_to_pes_11_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_63_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_63_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_63_io_to_pes_12_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_63_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_63_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_63_io_to_pes_13_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_63_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_63_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_63_io_to_pes_14_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_63_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_63_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_63_io_to_pes_15_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_63_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_63_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_63_io_to_pes_16_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_63_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_63_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_63_io_to_pes_17_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_63_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_63_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_63_io_to_pes_18_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_63_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_63_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_63_io_to_pes_19_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_63_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_63_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_63_io_to_pes_20_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_63_io_to_pes_21_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_63_io_to_pes_21_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_63_io_to_pes_21_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_63_io_to_mem_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_63_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_63_io_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_64_clock; // @[pe.scala 229:13]
  wire  PENetwork_64_reset; // @[pe.scala 229:13]
  wire  PENetwork_64_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_64_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_64_io_to_pes_0_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_64_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_64_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_64_io_to_pes_1_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_64_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_64_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_64_io_to_pes_2_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_64_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_64_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_64_io_to_pes_3_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_64_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_64_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_64_io_to_pes_4_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_64_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_64_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_64_io_to_pes_5_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_64_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_64_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_64_io_to_pes_6_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_64_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_64_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_64_io_to_pes_7_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_64_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_64_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_64_io_to_pes_8_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_64_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_64_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_64_io_to_pes_9_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_64_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_64_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_64_io_to_pes_10_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_64_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_64_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_64_io_to_pes_11_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_64_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_64_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_64_io_to_pes_12_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_64_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_64_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_64_io_to_pes_13_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_64_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_64_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_64_io_to_pes_14_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_64_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_64_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_64_io_to_pes_15_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_64_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_64_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_64_io_to_pes_16_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_64_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_64_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_64_io_to_pes_17_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_64_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_64_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_64_io_to_pes_18_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_64_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_64_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_64_io_to_pes_19_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_64_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_64_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_64_io_to_pes_20_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_64_io_to_pes_21_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_64_io_to_pes_21_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_64_io_to_pes_21_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_64_io_to_mem_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_64_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_64_io_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_65_clock; // @[pe.scala 229:13]
  wire  PENetwork_65_reset; // @[pe.scala 229:13]
  wire  PENetwork_65_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_65_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_65_io_to_pes_0_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_65_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_65_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_65_io_to_pes_1_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_65_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_65_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_65_io_to_pes_2_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_65_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_65_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_65_io_to_pes_3_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_65_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_65_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_65_io_to_pes_4_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_65_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_65_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_65_io_to_pes_5_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_65_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_65_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_65_io_to_pes_6_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_65_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_65_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_65_io_to_pes_7_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_65_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_65_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_65_io_to_pes_8_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_65_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_65_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_65_io_to_pes_9_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_65_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_65_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_65_io_to_pes_10_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_65_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_65_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_65_io_to_pes_11_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_65_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_65_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_65_io_to_pes_12_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_65_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_65_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_65_io_to_pes_13_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_65_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_65_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_65_io_to_pes_14_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_65_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_65_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_65_io_to_pes_15_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_65_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_65_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_65_io_to_pes_16_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_65_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_65_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_65_io_to_pes_17_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_65_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_65_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_65_io_to_pes_18_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_65_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_65_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_65_io_to_pes_19_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_65_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_65_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_65_io_to_pes_20_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_65_io_to_pes_21_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_65_io_to_pes_21_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_65_io_to_pes_21_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_65_io_to_mem_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_65_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_65_io_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_66_clock; // @[pe.scala 229:13]
  wire  PENetwork_66_reset; // @[pe.scala 229:13]
  wire  PENetwork_66_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_66_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_66_io_to_pes_0_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_66_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_66_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_66_io_to_pes_1_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_66_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_66_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_66_io_to_pes_2_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_66_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_66_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_66_io_to_pes_3_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_66_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_66_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_66_io_to_pes_4_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_66_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_66_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_66_io_to_pes_5_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_66_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_66_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_66_io_to_pes_6_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_66_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_66_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_66_io_to_pes_7_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_66_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_66_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_66_io_to_pes_8_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_66_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_66_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_66_io_to_pes_9_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_66_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_66_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_66_io_to_pes_10_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_66_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_66_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_66_io_to_pes_11_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_66_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_66_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_66_io_to_pes_12_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_66_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_66_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_66_io_to_pes_13_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_66_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_66_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_66_io_to_pes_14_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_66_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_66_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_66_io_to_pes_15_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_66_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_66_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_66_io_to_pes_16_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_66_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_66_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_66_io_to_pes_17_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_66_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_66_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_66_io_to_pes_18_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_66_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_66_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_66_io_to_pes_19_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_66_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_66_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_66_io_to_pes_20_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_66_io_to_pes_21_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_66_io_to_pes_21_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_66_io_to_pes_21_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_66_io_to_mem_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_66_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_66_io_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_67_clock; // @[pe.scala 229:13]
  wire  PENetwork_67_reset; // @[pe.scala 229:13]
  wire  PENetwork_67_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_67_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_67_io_to_pes_0_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_67_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_67_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_67_io_to_pes_1_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_67_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_67_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_67_io_to_pes_2_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_67_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_67_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_67_io_to_pes_3_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_67_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_67_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_67_io_to_pes_4_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_67_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_67_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_67_io_to_pes_5_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_67_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_67_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_67_io_to_pes_6_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_67_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_67_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_67_io_to_pes_7_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_67_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_67_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_67_io_to_pes_8_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_67_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_67_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_67_io_to_pes_9_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_67_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_67_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_67_io_to_pes_10_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_67_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_67_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_67_io_to_pes_11_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_67_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_67_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_67_io_to_pes_12_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_67_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_67_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_67_io_to_pes_13_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_67_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_67_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_67_io_to_pes_14_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_67_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_67_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_67_io_to_pes_15_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_67_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_67_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_67_io_to_pes_16_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_67_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_67_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_67_io_to_pes_17_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_67_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_67_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_67_io_to_pes_18_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_67_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_67_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_67_io_to_pes_19_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_67_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_67_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_67_io_to_pes_20_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_67_io_to_pes_21_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_67_io_to_pes_21_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_67_io_to_pes_21_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_67_io_to_mem_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_67_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_67_io_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_68_clock; // @[pe.scala 229:13]
  wire  PENetwork_68_reset; // @[pe.scala 229:13]
  wire  PENetwork_68_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_68_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_68_io_to_pes_0_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_68_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_68_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_68_io_to_pes_1_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_68_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_68_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_68_io_to_pes_2_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_68_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_68_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_68_io_to_pes_3_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_68_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_68_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_68_io_to_pes_4_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_68_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_68_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_68_io_to_pes_5_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_68_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_68_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_68_io_to_pes_6_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_68_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_68_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_68_io_to_pes_7_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_68_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_68_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_68_io_to_pes_8_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_68_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_68_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_68_io_to_pes_9_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_68_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_68_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_68_io_to_pes_10_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_68_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_68_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_68_io_to_pes_11_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_68_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_68_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_68_io_to_pes_12_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_68_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_68_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_68_io_to_pes_13_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_68_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_68_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_68_io_to_pes_14_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_68_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_68_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_68_io_to_pes_15_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_68_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_68_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_68_io_to_pes_16_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_68_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_68_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_68_io_to_pes_17_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_68_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_68_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_68_io_to_pes_18_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_68_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_68_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_68_io_to_pes_19_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_68_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_68_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_68_io_to_pes_20_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_68_io_to_pes_21_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_68_io_to_pes_21_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_68_io_to_pes_21_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_68_io_to_mem_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_68_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_68_io_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_69_clock; // @[pe.scala 229:13]
  wire  PENetwork_69_reset; // @[pe.scala 229:13]
  wire  PENetwork_69_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_69_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_69_io_to_pes_0_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_69_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_69_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_69_io_to_pes_1_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_69_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_69_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_69_io_to_pes_2_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_69_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_69_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_69_io_to_pes_3_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_69_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_69_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_69_io_to_pes_4_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_69_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_69_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_69_io_to_pes_5_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_69_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_69_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_69_io_to_pes_6_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_69_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_69_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_69_io_to_pes_7_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_69_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_69_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_69_io_to_pes_8_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_69_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_69_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_69_io_to_pes_9_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_69_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_69_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_69_io_to_pes_10_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_69_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_69_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_69_io_to_pes_11_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_69_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_69_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_69_io_to_pes_12_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_69_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_69_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_69_io_to_pes_13_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_69_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_69_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_69_io_to_pes_14_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_69_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_69_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_69_io_to_pes_15_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_69_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_69_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_69_io_to_pes_16_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_69_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_69_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_69_io_to_pes_17_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_69_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_69_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_69_io_to_pes_18_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_69_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_69_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_69_io_to_pes_19_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_69_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_69_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_69_io_to_pes_20_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_69_io_to_pes_21_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_69_io_to_pes_21_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_69_io_to_pes_21_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_69_io_to_mem_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_69_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_69_io_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_70_clock; // @[pe.scala 229:13]
  wire  PENetwork_70_reset; // @[pe.scala 229:13]
  wire  PENetwork_70_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_70_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_70_io_to_pes_0_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_70_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_70_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_70_io_to_pes_1_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_70_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_70_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_70_io_to_pes_2_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_70_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_70_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_70_io_to_pes_3_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_70_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_70_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_70_io_to_pes_4_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_70_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_70_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_70_io_to_pes_5_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_70_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_70_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_70_io_to_pes_6_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_70_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_70_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_70_io_to_pes_7_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_70_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_70_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_70_io_to_pes_8_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_70_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_70_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_70_io_to_pes_9_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_70_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_70_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_70_io_to_pes_10_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_70_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_70_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_70_io_to_pes_11_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_70_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_70_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_70_io_to_pes_12_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_70_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_70_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_70_io_to_pes_13_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_70_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_70_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_70_io_to_pes_14_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_70_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_70_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_70_io_to_pes_15_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_70_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_70_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_70_io_to_pes_16_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_70_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_70_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_70_io_to_pes_17_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_70_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_70_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_70_io_to_pes_18_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_70_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_70_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_70_io_to_pes_19_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_70_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_70_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_70_io_to_pes_20_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_70_io_to_pes_21_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_70_io_to_pes_21_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_70_io_to_pes_21_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_70_io_to_mem_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_70_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_70_io_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_71_clock; // @[pe.scala 229:13]
  wire  PENetwork_71_reset; // @[pe.scala 229:13]
  wire  PENetwork_71_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_71_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_71_io_to_pes_0_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_71_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_71_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_71_io_to_pes_1_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_71_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_71_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_71_io_to_pes_2_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_71_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_71_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_71_io_to_pes_3_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_71_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_71_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_71_io_to_pes_4_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_71_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_71_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_71_io_to_pes_5_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_71_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_71_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_71_io_to_pes_6_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_71_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_71_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_71_io_to_pes_7_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_71_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_71_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_71_io_to_pes_8_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_71_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_71_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_71_io_to_pes_9_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_71_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_71_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_71_io_to_pes_10_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_71_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_71_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_71_io_to_pes_11_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_71_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_71_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_71_io_to_pes_12_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_71_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_71_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_71_io_to_pes_13_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_71_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_71_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_71_io_to_pes_14_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_71_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_71_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_71_io_to_pes_15_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_71_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_71_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_71_io_to_pes_16_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_71_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_71_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_71_io_to_pes_17_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_71_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_71_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_71_io_to_pes_18_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_71_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_71_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_71_io_to_pes_19_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_71_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_71_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_71_io_to_pes_20_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_71_io_to_pes_21_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_71_io_to_pes_21_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_71_io_to_pes_21_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_71_io_to_mem_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_71_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_71_io_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_72_clock; // @[pe.scala 229:13]
  wire  PENetwork_72_reset; // @[pe.scala 229:13]
  wire  PENetwork_72_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_72_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_72_io_to_pes_0_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_72_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_72_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_72_io_to_pes_1_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_72_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_72_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_72_io_to_pes_2_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_72_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_72_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_72_io_to_pes_3_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_72_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_72_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_72_io_to_pes_4_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_72_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_72_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_72_io_to_pes_5_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_72_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_72_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_72_io_to_pes_6_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_72_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_72_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_72_io_to_pes_7_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_72_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_72_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_72_io_to_pes_8_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_72_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_72_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_72_io_to_pes_9_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_72_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_72_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_72_io_to_pes_10_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_72_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_72_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_72_io_to_pes_11_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_72_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_72_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_72_io_to_pes_12_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_72_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_72_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_72_io_to_pes_13_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_72_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_72_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_72_io_to_pes_14_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_72_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_72_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_72_io_to_pes_15_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_72_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_72_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_72_io_to_pes_16_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_72_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_72_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_72_io_to_pes_17_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_72_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_72_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_72_io_to_pes_18_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_72_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_72_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_72_io_to_pes_19_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_72_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_72_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_72_io_to_pes_20_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_72_io_to_pes_21_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_72_io_to_pes_21_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_72_io_to_pes_21_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_72_io_to_mem_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_72_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_72_io_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_73_clock; // @[pe.scala 229:13]
  wire  PENetwork_73_reset; // @[pe.scala 229:13]
  wire  PENetwork_73_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_73_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_73_io_to_pes_0_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_73_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_73_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_73_io_to_pes_1_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_73_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_73_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_73_io_to_pes_2_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_73_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_73_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_73_io_to_pes_3_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_73_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_73_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_73_io_to_pes_4_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_73_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_73_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_73_io_to_pes_5_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_73_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_73_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_73_io_to_pes_6_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_73_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_73_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_73_io_to_pes_7_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_73_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_73_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_73_io_to_pes_8_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_73_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_73_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_73_io_to_pes_9_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_73_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_73_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_73_io_to_pes_10_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_73_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_73_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_73_io_to_pes_11_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_73_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_73_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_73_io_to_pes_12_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_73_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_73_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_73_io_to_pes_13_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_73_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_73_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_73_io_to_pes_14_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_73_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_73_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_73_io_to_pes_15_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_73_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_73_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_73_io_to_pes_16_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_73_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_73_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_73_io_to_pes_17_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_73_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_73_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_73_io_to_pes_18_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_73_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_73_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_73_io_to_pes_19_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_73_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_73_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_73_io_to_pes_20_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_73_io_to_pes_21_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_73_io_to_pes_21_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_73_io_to_pes_21_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_73_io_to_mem_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_73_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_73_io_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_74_clock; // @[pe.scala 229:13]
  wire  PENetwork_74_reset; // @[pe.scala 229:13]
  wire  PENetwork_74_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_74_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_74_io_to_pes_0_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_74_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_74_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_74_io_to_pes_1_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_74_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_74_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_74_io_to_pes_2_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_74_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_74_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_74_io_to_pes_3_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_74_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_74_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_74_io_to_pes_4_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_74_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_74_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_74_io_to_pes_5_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_74_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_74_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_74_io_to_pes_6_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_74_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_74_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_74_io_to_pes_7_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_74_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_74_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_74_io_to_pes_8_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_74_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_74_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_74_io_to_pes_9_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_74_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_74_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_74_io_to_pes_10_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_74_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_74_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_74_io_to_pes_11_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_74_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_74_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_74_io_to_pes_12_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_74_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_74_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_74_io_to_pes_13_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_74_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_74_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_74_io_to_pes_14_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_74_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_74_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_74_io_to_pes_15_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_74_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_74_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_74_io_to_pes_16_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_74_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_74_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_74_io_to_pes_17_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_74_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_74_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_74_io_to_pes_18_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_74_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_74_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_74_io_to_pes_19_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_74_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_74_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_74_io_to_pes_20_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_74_io_to_pes_21_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_74_io_to_pes_21_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_74_io_to_pes_21_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_74_io_to_mem_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_74_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_74_io_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_75_clock; // @[pe.scala 229:13]
  wire  PENetwork_75_reset; // @[pe.scala 229:13]
  wire  PENetwork_75_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_75_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_75_io_to_pes_0_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_75_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_75_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_75_io_to_pes_1_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_75_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_75_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_75_io_to_pes_2_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_75_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_75_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_75_io_to_pes_3_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_75_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_75_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_75_io_to_pes_4_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_75_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_75_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_75_io_to_pes_5_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_75_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_75_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_75_io_to_pes_6_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_75_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_75_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_75_io_to_pes_7_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_75_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_75_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_75_io_to_pes_8_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_75_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_75_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_75_io_to_pes_9_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_75_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_75_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_75_io_to_pes_10_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_75_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_75_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_75_io_to_pes_11_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_75_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_75_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_75_io_to_pes_12_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_75_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_75_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_75_io_to_pes_13_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_75_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_75_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_75_io_to_pes_14_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_75_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_75_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_75_io_to_pes_15_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_75_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_75_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_75_io_to_pes_16_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_75_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_75_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_75_io_to_pes_17_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_75_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_75_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_75_io_to_pes_18_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_75_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_75_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_75_io_to_pes_19_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_75_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_75_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_75_io_to_pes_20_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_75_io_to_pes_21_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_75_io_to_pes_21_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_75_io_to_pes_21_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_75_io_to_mem_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_75_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_75_io_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_76_clock; // @[pe.scala 229:13]
  wire  PENetwork_76_reset; // @[pe.scala 229:13]
  wire  PENetwork_76_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_76_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_76_io_to_pes_0_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_76_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_76_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_76_io_to_pes_1_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_76_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_76_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_76_io_to_pes_2_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_76_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_76_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_76_io_to_pes_3_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_76_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_76_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_76_io_to_pes_4_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_76_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_76_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_76_io_to_pes_5_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_76_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_76_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_76_io_to_pes_6_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_76_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_76_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_76_io_to_pes_7_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_76_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_76_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_76_io_to_pes_8_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_76_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_76_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_76_io_to_pes_9_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_76_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_76_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_76_io_to_pes_10_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_76_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_76_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_76_io_to_pes_11_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_76_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_76_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_76_io_to_pes_12_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_76_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_76_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_76_io_to_pes_13_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_76_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_76_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_76_io_to_pes_14_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_76_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_76_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_76_io_to_pes_15_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_76_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_76_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_76_io_to_pes_16_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_76_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_76_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_76_io_to_pes_17_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_76_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_76_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_76_io_to_pes_18_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_76_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_76_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_76_io_to_pes_19_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_76_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_76_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_76_io_to_pes_20_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_76_io_to_pes_21_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_76_io_to_pes_21_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_76_io_to_pes_21_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_76_io_to_mem_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_76_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_76_io_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_77_clock; // @[pe.scala 229:13]
  wire  PENetwork_77_reset; // @[pe.scala 229:13]
  wire  PENetwork_77_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_77_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_77_io_to_pes_0_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_77_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_77_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_77_io_to_pes_1_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_77_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_77_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_77_io_to_pes_2_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_77_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_77_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_77_io_to_pes_3_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_77_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_77_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_77_io_to_pes_4_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_77_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_77_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_77_io_to_pes_5_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_77_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_77_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_77_io_to_pes_6_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_77_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_77_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_77_io_to_pes_7_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_77_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_77_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_77_io_to_pes_8_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_77_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_77_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_77_io_to_pes_9_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_77_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_77_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_77_io_to_pes_10_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_77_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_77_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_77_io_to_pes_11_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_77_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_77_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_77_io_to_pes_12_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_77_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_77_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_77_io_to_pes_13_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_77_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_77_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_77_io_to_pes_14_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_77_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_77_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_77_io_to_pes_15_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_77_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_77_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_77_io_to_pes_16_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_77_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_77_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_77_io_to_pes_17_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_77_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_77_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_77_io_to_pes_18_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_77_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_77_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_77_io_to_pes_19_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_77_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_77_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_77_io_to_pes_20_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_77_io_to_pes_21_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_77_io_to_pes_21_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_77_io_to_pes_21_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_77_io_to_mem_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_77_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_77_io_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_78_clock; // @[pe.scala 229:13]
  wire  PENetwork_78_reset; // @[pe.scala 229:13]
  wire  PENetwork_78_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_78_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_78_io_to_pes_0_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_78_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_78_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_78_io_to_pes_1_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_78_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_78_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_78_io_to_pes_2_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_78_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_78_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_78_io_to_pes_3_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_78_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_78_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_78_io_to_pes_4_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_78_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_78_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_78_io_to_pes_5_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_78_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_78_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_78_io_to_pes_6_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_78_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_78_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_78_io_to_pes_7_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_78_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_78_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_78_io_to_pes_8_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_78_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_78_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_78_io_to_pes_9_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_78_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_78_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_78_io_to_pes_10_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_78_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_78_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_78_io_to_pes_11_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_78_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_78_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_78_io_to_pes_12_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_78_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_78_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_78_io_to_pes_13_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_78_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_78_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_78_io_to_pes_14_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_78_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_78_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_78_io_to_pes_15_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_78_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_78_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_78_io_to_pes_16_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_78_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_78_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_78_io_to_pes_17_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_78_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_78_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_78_io_to_pes_18_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_78_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_78_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_78_io_to_pes_19_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_78_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_78_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_78_io_to_pes_20_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_78_io_to_pes_21_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_78_io_to_pes_21_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_78_io_to_pes_21_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_78_io_to_mem_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_78_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_78_io_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_79_clock; // @[pe.scala 229:13]
  wire  PENetwork_79_reset; // @[pe.scala 229:13]
  wire  PENetwork_79_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_79_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_79_io_to_pes_0_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_79_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_79_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_79_io_to_pes_1_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_79_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_79_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_79_io_to_pes_2_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_79_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_79_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_79_io_to_pes_3_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_79_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_79_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_79_io_to_pes_4_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_79_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_79_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_79_io_to_pes_5_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_79_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_79_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_79_io_to_pes_6_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_79_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_79_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_79_io_to_pes_7_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_79_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_79_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_79_io_to_pes_8_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_79_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_79_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_79_io_to_pes_9_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_79_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_79_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_79_io_to_pes_10_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_79_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_79_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_79_io_to_pes_11_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_79_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_79_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_79_io_to_pes_12_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_79_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_79_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_79_io_to_pes_13_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_79_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_79_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_79_io_to_pes_14_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_79_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_79_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_79_io_to_pes_15_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_79_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_79_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_79_io_to_pes_16_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_79_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_79_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_79_io_to_pes_17_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_79_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_79_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_79_io_to_pes_18_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_79_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_79_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_79_io_to_pes_19_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_79_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_79_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_79_io_to_pes_20_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_79_io_to_pes_21_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_79_io_to_pes_21_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_79_io_to_pes_21_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_79_io_to_mem_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_79_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_79_io_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_80_clock; // @[pe.scala 229:13]
  wire  PENetwork_80_reset; // @[pe.scala 229:13]
  wire  PENetwork_80_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_80_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_80_io_to_pes_0_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_80_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_80_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_80_io_to_pes_1_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_80_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_80_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_80_io_to_pes_2_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_80_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_80_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_80_io_to_pes_3_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_80_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_80_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_80_io_to_pes_4_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_80_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_80_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_80_io_to_pes_5_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_80_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_80_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_80_io_to_pes_6_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_80_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_80_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_80_io_to_pes_7_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_80_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_80_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_80_io_to_pes_8_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_80_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_80_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_80_io_to_pes_9_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_80_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_80_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_80_io_to_pes_10_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_80_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_80_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_80_io_to_pes_11_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_80_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_80_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_80_io_to_pes_12_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_80_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_80_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_80_io_to_pes_13_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_80_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_80_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_80_io_to_pes_14_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_80_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_80_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_80_io_to_pes_15_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_80_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_80_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_80_io_to_pes_16_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_80_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_80_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_80_io_to_pes_17_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_80_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_80_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_80_io_to_pes_18_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_80_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_80_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_80_io_to_pes_19_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_80_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_80_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_80_io_to_pes_20_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_80_io_to_pes_21_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_80_io_to_pes_21_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_80_io_to_pes_21_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_80_io_to_mem_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_80_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_80_io_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_81_clock; // @[pe.scala 229:13]
  wire  PENetwork_81_reset; // @[pe.scala 229:13]
  wire  PENetwork_81_io_to_pes_0_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_81_io_to_pes_0_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_81_io_to_pes_0_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_81_io_to_pes_1_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_81_io_to_pes_1_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_81_io_to_pes_1_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_81_io_to_pes_2_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_81_io_to_pes_2_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_81_io_to_pes_2_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_81_io_to_pes_3_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_81_io_to_pes_3_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_81_io_to_pes_3_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_81_io_to_pes_4_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_81_io_to_pes_4_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_81_io_to_pes_4_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_81_io_to_pes_5_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_81_io_to_pes_5_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_81_io_to_pes_5_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_81_io_to_pes_6_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_81_io_to_pes_6_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_81_io_to_pes_6_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_81_io_to_pes_7_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_81_io_to_pes_7_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_81_io_to_pes_7_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_81_io_to_pes_8_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_81_io_to_pes_8_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_81_io_to_pes_8_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_81_io_to_pes_9_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_81_io_to_pes_9_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_81_io_to_pes_9_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_81_io_to_pes_10_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_81_io_to_pes_10_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_81_io_to_pes_10_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_81_io_to_pes_11_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_81_io_to_pes_11_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_81_io_to_pes_11_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_81_io_to_pes_12_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_81_io_to_pes_12_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_81_io_to_pes_12_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_81_io_to_pes_13_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_81_io_to_pes_13_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_81_io_to_pes_13_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_81_io_to_pes_14_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_81_io_to_pes_14_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_81_io_to_pes_14_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_81_io_to_pes_15_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_81_io_to_pes_15_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_81_io_to_pes_15_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_81_io_to_pes_16_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_81_io_to_pes_16_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_81_io_to_pes_16_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_81_io_to_pes_17_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_81_io_to_pes_17_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_81_io_to_pes_17_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_81_io_to_pes_18_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_81_io_to_pes_18_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_81_io_to_pes_18_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_81_io_to_pes_19_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_81_io_to_pes_19_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_81_io_to_pes_19_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_81_io_to_pes_20_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_81_io_to_pes_20_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_81_io_to_pes_20_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_81_io_to_pes_21_out_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_81_io_to_pes_21_out_bits; // @[pe.scala 229:13]
  wire  PENetwork_81_io_to_pes_21_sig_stat2trans; // @[pe.scala 229:13]
  wire  PENetwork_81_io_to_mem_valid; // @[pe.scala 229:13]
  wire [127:0] PENetwork_81_io_to_mem_bits; // @[pe.scala 229:13]
  wire  PENetwork_81_io_sig_stat2trans; // @[pe.scala 229:13]
  wire  MemController_clock; // @[pe.scala 303:15]
  wire  MemController_reset; // @[pe.scala 303:15]
  wire  MemController_io_rd_valid; // @[pe.scala 303:15]
  wire  MemController_io_wr_valid; // @[pe.scala 303:15]
  wire  MemController_io_rd_data_valid; // @[pe.scala 303:15]
  wire [15:0] MemController_io_rd_data_bits; // @[pe.scala 303:15]
  wire  MemController_io_wr_data_valid; // @[pe.scala 303:15]
  wire [15:0] MemController_io_wr_data_bits; // @[pe.scala 303:15]
  wire  MemController_1_clock; // @[pe.scala 303:15]
  wire  MemController_1_reset; // @[pe.scala 303:15]
  wire  MemController_1_io_rd_valid; // @[pe.scala 303:15]
  wire  MemController_1_io_wr_valid; // @[pe.scala 303:15]
  wire  MemController_1_io_rd_data_valid; // @[pe.scala 303:15]
  wire [15:0] MemController_1_io_rd_data_bits; // @[pe.scala 303:15]
  wire  MemController_1_io_wr_data_valid; // @[pe.scala 303:15]
  wire [15:0] MemController_1_io_wr_data_bits; // @[pe.scala 303:15]
  wire  MemController_2_clock; // @[pe.scala 303:15]
  wire  MemController_2_reset; // @[pe.scala 303:15]
  wire  MemController_2_io_rd_valid; // @[pe.scala 303:15]
  wire  MemController_2_io_wr_valid; // @[pe.scala 303:15]
  wire  MemController_2_io_rd_data_valid; // @[pe.scala 303:15]
  wire [15:0] MemController_2_io_rd_data_bits; // @[pe.scala 303:15]
  wire  MemController_2_io_wr_data_valid; // @[pe.scala 303:15]
  wire [15:0] MemController_2_io_wr_data_bits; // @[pe.scala 303:15]
  wire  MemController_3_clock; // @[pe.scala 303:15]
  wire  MemController_3_reset; // @[pe.scala 303:15]
  wire  MemController_3_io_rd_valid; // @[pe.scala 303:15]
  wire  MemController_3_io_wr_valid; // @[pe.scala 303:15]
  wire  MemController_3_io_rd_data_valid; // @[pe.scala 303:15]
  wire [15:0] MemController_3_io_rd_data_bits; // @[pe.scala 303:15]
  wire  MemController_3_io_wr_data_valid; // @[pe.scala 303:15]
  wire [15:0] MemController_3_io_wr_data_bits; // @[pe.scala 303:15]
  wire  MemController_4_clock; // @[pe.scala 303:15]
  wire  MemController_4_reset; // @[pe.scala 303:15]
  wire  MemController_4_io_rd_valid; // @[pe.scala 303:15]
  wire  MemController_4_io_wr_valid; // @[pe.scala 303:15]
  wire  MemController_4_io_rd_data_valid; // @[pe.scala 303:15]
  wire [15:0] MemController_4_io_rd_data_bits; // @[pe.scala 303:15]
  wire  MemController_4_io_wr_data_valid; // @[pe.scala 303:15]
  wire [15:0] MemController_4_io_wr_data_bits; // @[pe.scala 303:15]
  wire  MemController_5_clock; // @[pe.scala 303:15]
  wire  MemController_5_reset; // @[pe.scala 303:15]
  wire  MemController_5_io_rd_valid; // @[pe.scala 303:15]
  wire  MemController_5_io_wr_valid; // @[pe.scala 303:15]
  wire  MemController_5_io_rd_data_valid; // @[pe.scala 303:15]
  wire [15:0] MemController_5_io_rd_data_bits; // @[pe.scala 303:15]
  wire  MemController_5_io_wr_data_valid; // @[pe.scala 303:15]
  wire [15:0] MemController_5_io_wr_data_bits; // @[pe.scala 303:15]
  wire  MemController_6_clock; // @[pe.scala 303:15]
  wire  MemController_6_reset; // @[pe.scala 303:15]
  wire  MemController_6_io_rd_valid; // @[pe.scala 303:15]
  wire  MemController_6_io_wr_valid; // @[pe.scala 303:15]
  wire  MemController_6_io_rd_data_valid; // @[pe.scala 303:15]
  wire [15:0] MemController_6_io_rd_data_bits; // @[pe.scala 303:15]
  wire  MemController_6_io_wr_data_valid; // @[pe.scala 303:15]
  wire [15:0] MemController_6_io_wr_data_bits; // @[pe.scala 303:15]
  wire  MemController_7_clock; // @[pe.scala 303:15]
  wire  MemController_7_reset; // @[pe.scala 303:15]
  wire  MemController_7_io_rd_valid; // @[pe.scala 303:15]
  wire  MemController_7_io_wr_valid; // @[pe.scala 303:15]
  wire  MemController_7_io_rd_data_valid; // @[pe.scala 303:15]
  wire [15:0] MemController_7_io_rd_data_bits; // @[pe.scala 303:15]
  wire  MemController_7_io_wr_data_valid; // @[pe.scala 303:15]
  wire [15:0] MemController_7_io_wr_data_bits; // @[pe.scala 303:15]
  wire  MemController_8_clock; // @[pe.scala 303:15]
  wire  MemController_8_reset; // @[pe.scala 303:15]
  wire  MemController_8_io_rd_valid; // @[pe.scala 303:15]
  wire  MemController_8_io_wr_valid; // @[pe.scala 303:15]
  wire  MemController_8_io_rd_data_valid; // @[pe.scala 303:15]
  wire [15:0] MemController_8_io_rd_data_bits; // @[pe.scala 303:15]
  wire  MemController_8_io_wr_data_valid; // @[pe.scala 303:15]
  wire [15:0] MemController_8_io_wr_data_bits; // @[pe.scala 303:15]
  wire  MemController_9_clock; // @[pe.scala 303:15]
  wire  MemController_9_reset; // @[pe.scala 303:15]
  wire  MemController_9_io_rd_valid; // @[pe.scala 303:15]
  wire  MemController_9_io_wr_valid; // @[pe.scala 303:15]
  wire  MemController_9_io_rd_data_valid; // @[pe.scala 303:15]
  wire [15:0] MemController_9_io_rd_data_bits; // @[pe.scala 303:15]
  wire  MemController_9_io_wr_data_valid; // @[pe.scala 303:15]
  wire [15:0] MemController_9_io_wr_data_bits; // @[pe.scala 303:15]
  wire  MemController_10_clock; // @[pe.scala 303:15]
  wire  MemController_10_reset; // @[pe.scala 303:15]
  wire  MemController_10_io_rd_valid; // @[pe.scala 303:15]
  wire  MemController_10_io_wr_valid; // @[pe.scala 303:15]
  wire  MemController_10_io_rd_data_valid; // @[pe.scala 303:15]
  wire [15:0] MemController_10_io_rd_data_bits; // @[pe.scala 303:15]
  wire  MemController_10_io_wr_data_valid; // @[pe.scala 303:15]
  wire [15:0] MemController_10_io_wr_data_bits; // @[pe.scala 303:15]
  wire  MemController_11_clock; // @[pe.scala 303:15]
  wire  MemController_11_reset; // @[pe.scala 303:15]
  wire  MemController_11_io_rd_valid; // @[pe.scala 303:15]
  wire  MemController_11_io_wr_valid; // @[pe.scala 303:15]
  wire  MemController_11_io_rd_data_valid; // @[pe.scala 303:15]
  wire [15:0] MemController_11_io_rd_data_bits; // @[pe.scala 303:15]
  wire  MemController_11_io_wr_data_valid; // @[pe.scala 303:15]
  wire [15:0] MemController_11_io_wr_data_bits; // @[pe.scala 303:15]
  wire  MemController_12_clock; // @[pe.scala 303:15]
  wire  MemController_12_reset; // @[pe.scala 303:15]
  wire  MemController_12_io_rd_valid; // @[pe.scala 303:15]
  wire  MemController_12_io_wr_valid; // @[pe.scala 303:15]
  wire  MemController_12_io_rd_data_valid; // @[pe.scala 303:15]
  wire [15:0] MemController_12_io_rd_data_bits; // @[pe.scala 303:15]
  wire  MemController_12_io_wr_data_valid; // @[pe.scala 303:15]
  wire [15:0] MemController_12_io_wr_data_bits; // @[pe.scala 303:15]
  wire  MemController_13_clock; // @[pe.scala 303:15]
  wire  MemController_13_reset; // @[pe.scala 303:15]
  wire  MemController_13_io_rd_valid; // @[pe.scala 303:15]
  wire  MemController_13_io_wr_valid; // @[pe.scala 303:15]
  wire  MemController_13_io_rd_data_valid; // @[pe.scala 303:15]
  wire [15:0] MemController_13_io_rd_data_bits; // @[pe.scala 303:15]
  wire  MemController_13_io_wr_data_valid; // @[pe.scala 303:15]
  wire [15:0] MemController_13_io_wr_data_bits; // @[pe.scala 303:15]
  wire  MemController_14_clock; // @[pe.scala 303:15]
  wire  MemController_14_reset; // @[pe.scala 303:15]
  wire  MemController_14_io_rd_valid; // @[pe.scala 303:15]
  wire  MemController_14_io_wr_valid; // @[pe.scala 303:15]
  wire  MemController_14_io_rd_data_valid; // @[pe.scala 303:15]
  wire [15:0] MemController_14_io_rd_data_bits; // @[pe.scala 303:15]
  wire  MemController_14_io_wr_data_valid; // @[pe.scala 303:15]
  wire [15:0] MemController_14_io_wr_data_bits; // @[pe.scala 303:15]
  wire  MemController_15_clock; // @[pe.scala 303:15]
  wire  MemController_15_reset; // @[pe.scala 303:15]
  wire  MemController_15_io_rd_valid; // @[pe.scala 303:15]
  wire  MemController_15_io_wr_valid; // @[pe.scala 303:15]
  wire  MemController_15_io_rd_data_valid; // @[pe.scala 303:15]
  wire [15:0] MemController_15_io_rd_data_bits; // @[pe.scala 303:15]
  wire  MemController_15_io_wr_data_valid; // @[pe.scala 303:15]
  wire [15:0] MemController_15_io_wr_data_bits; // @[pe.scala 303:15]
  wire  MemController_16_clock; // @[pe.scala 303:15]
  wire  MemController_16_reset; // @[pe.scala 303:15]
  wire  MemController_16_io_rd_valid; // @[pe.scala 303:15]
  wire  MemController_16_io_wr_valid; // @[pe.scala 303:15]
  wire  MemController_16_io_rd_data_valid; // @[pe.scala 303:15]
  wire [15:0] MemController_16_io_rd_data_bits; // @[pe.scala 303:15]
  wire  MemController_16_io_wr_data_valid; // @[pe.scala 303:15]
  wire [15:0] MemController_16_io_wr_data_bits; // @[pe.scala 303:15]
  wire  MemController_17_clock; // @[pe.scala 303:15]
  wire  MemController_17_reset; // @[pe.scala 303:15]
  wire  MemController_17_io_rd_valid; // @[pe.scala 303:15]
  wire  MemController_17_io_wr_valid; // @[pe.scala 303:15]
  wire  MemController_17_io_rd_data_valid; // @[pe.scala 303:15]
  wire [15:0] MemController_17_io_rd_data_bits; // @[pe.scala 303:15]
  wire  MemController_17_io_wr_data_valid; // @[pe.scala 303:15]
  wire [15:0] MemController_17_io_wr_data_bits; // @[pe.scala 303:15]
  wire  MemController_18_clock; // @[pe.scala 303:15]
  wire  MemController_18_reset; // @[pe.scala 303:15]
  wire  MemController_18_io_rd_valid; // @[pe.scala 303:15]
  wire  MemController_18_io_wr_valid; // @[pe.scala 303:15]
  wire  MemController_18_io_rd_data_valid; // @[pe.scala 303:15]
  wire [15:0] MemController_18_io_rd_data_bits; // @[pe.scala 303:15]
  wire  MemController_18_io_wr_data_valid; // @[pe.scala 303:15]
  wire [15:0] MemController_18_io_wr_data_bits; // @[pe.scala 303:15]
  wire  MemController_19_clock; // @[pe.scala 303:15]
  wire  MemController_19_reset; // @[pe.scala 303:15]
  wire  MemController_19_io_rd_valid; // @[pe.scala 303:15]
  wire  MemController_19_io_wr_valid; // @[pe.scala 303:15]
  wire  MemController_19_io_rd_data_valid; // @[pe.scala 303:15]
  wire [15:0] MemController_19_io_rd_data_bits; // @[pe.scala 303:15]
  wire  MemController_19_io_wr_data_valid; // @[pe.scala 303:15]
  wire [15:0] MemController_19_io_wr_data_bits; // @[pe.scala 303:15]
  wire  MemController_20_clock; // @[pe.scala 303:15]
  wire  MemController_20_reset; // @[pe.scala 303:15]
  wire  MemController_20_io_rd_valid; // @[pe.scala 303:15]
  wire  MemController_20_io_wr_valid; // @[pe.scala 303:15]
  wire  MemController_20_io_rd_data_valid; // @[pe.scala 303:15]
  wire [15:0] MemController_20_io_rd_data_bits; // @[pe.scala 303:15]
  wire  MemController_20_io_wr_data_valid; // @[pe.scala 303:15]
  wire [15:0] MemController_20_io_wr_data_bits; // @[pe.scala 303:15]
  wire  MemController_21_clock; // @[pe.scala 303:15]
  wire  MemController_21_reset; // @[pe.scala 303:15]
  wire  MemController_21_io_rd_valid; // @[pe.scala 303:15]
  wire  MemController_21_io_wr_valid; // @[pe.scala 303:15]
  wire  MemController_21_io_rd_data_valid; // @[pe.scala 303:15]
  wire [15:0] MemController_21_io_rd_data_bits; // @[pe.scala 303:15]
  wire  MemController_21_io_wr_data_valid; // @[pe.scala 303:15]
  wire [15:0] MemController_21_io_wr_data_bits; // @[pe.scala 303:15]
  wire  MemController_22_clock; // @[pe.scala 303:15]
  wire  MemController_22_reset; // @[pe.scala 303:15]
  wire  MemController_22_io_rd_valid; // @[pe.scala 303:15]
  wire  MemController_22_io_wr_valid; // @[pe.scala 303:15]
  wire  MemController_22_io_rd_data_valid; // @[pe.scala 303:15]
  wire [127:0] MemController_22_io_rd_data_bits; // @[pe.scala 303:15]
  wire  MemController_22_io_wr_data_valid; // @[pe.scala 303:15]
  wire [127:0] MemController_22_io_wr_data_bits; // @[pe.scala 303:15]
  wire  MemController_23_clock; // @[pe.scala 303:15]
  wire  MemController_23_reset; // @[pe.scala 303:15]
  wire  MemController_23_io_rd_valid; // @[pe.scala 303:15]
  wire  MemController_23_io_wr_valid; // @[pe.scala 303:15]
  wire  MemController_23_io_rd_data_valid; // @[pe.scala 303:15]
  wire [127:0] MemController_23_io_rd_data_bits; // @[pe.scala 303:15]
  wire  MemController_23_io_wr_data_valid; // @[pe.scala 303:15]
  wire [127:0] MemController_23_io_wr_data_bits; // @[pe.scala 303:15]
  wire  MemController_24_clock; // @[pe.scala 303:15]
  wire  MemController_24_reset; // @[pe.scala 303:15]
  wire  MemController_24_io_rd_valid; // @[pe.scala 303:15]
  wire  MemController_24_io_wr_valid; // @[pe.scala 303:15]
  wire  MemController_24_io_rd_data_valid; // @[pe.scala 303:15]
  wire [127:0] MemController_24_io_rd_data_bits; // @[pe.scala 303:15]
  wire  MemController_24_io_wr_data_valid; // @[pe.scala 303:15]
  wire [127:0] MemController_24_io_wr_data_bits; // @[pe.scala 303:15]
  wire  MemController_25_clock; // @[pe.scala 303:15]
  wire  MemController_25_reset; // @[pe.scala 303:15]
  wire  MemController_25_io_rd_valid; // @[pe.scala 303:15]
  wire  MemController_25_io_wr_valid; // @[pe.scala 303:15]
  wire  MemController_25_io_rd_data_valid; // @[pe.scala 303:15]
  wire [127:0] MemController_25_io_rd_data_bits; // @[pe.scala 303:15]
  wire  MemController_25_io_wr_data_valid; // @[pe.scala 303:15]
  wire [127:0] MemController_25_io_wr_data_bits; // @[pe.scala 303:15]
  wire  MemController_26_clock; // @[pe.scala 303:15]
  wire  MemController_26_reset; // @[pe.scala 303:15]
  wire  MemController_26_io_rd_valid; // @[pe.scala 303:15]
  wire  MemController_26_io_wr_valid; // @[pe.scala 303:15]
  wire  MemController_26_io_rd_data_valid; // @[pe.scala 303:15]
  wire [127:0] MemController_26_io_rd_data_bits; // @[pe.scala 303:15]
  wire  MemController_26_io_wr_data_valid; // @[pe.scala 303:15]
  wire [127:0] MemController_26_io_wr_data_bits; // @[pe.scala 303:15]
  wire  MemController_27_clock; // @[pe.scala 303:15]
  wire  MemController_27_reset; // @[pe.scala 303:15]
  wire  MemController_27_io_rd_valid; // @[pe.scala 303:15]
  wire  MemController_27_io_wr_valid; // @[pe.scala 303:15]
  wire  MemController_27_io_rd_data_valid; // @[pe.scala 303:15]
  wire [127:0] MemController_27_io_rd_data_bits; // @[pe.scala 303:15]
  wire  MemController_27_io_wr_data_valid; // @[pe.scala 303:15]
  wire [127:0] MemController_27_io_wr_data_bits; // @[pe.scala 303:15]
  wire  MemController_28_clock; // @[pe.scala 303:15]
  wire  MemController_28_reset; // @[pe.scala 303:15]
  wire  MemController_28_io_rd_valid; // @[pe.scala 303:15]
  wire  MemController_28_io_wr_valid; // @[pe.scala 303:15]
  wire  MemController_28_io_rd_data_valid; // @[pe.scala 303:15]
  wire [127:0] MemController_28_io_rd_data_bits; // @[pe.scala 303:15]
  wire  MemController_28_io_wr_data_valid; // @[pe.scala 303:15]
  wire [127:0] MemController_28_io_wr_data_bits; // @[pe.scala 303:15]
  wire  MemController_29_clock; // @[pe.scala 303:15]
  wire  MemController_29_reset; // @[pe.scala 303:15]
  wire  MemController_29_io_rd_valid; // @[pe.scala 303:15]
  wire  MemController_29_io_wr_valid; // @[pe.scala 303:15]
  wire  MemController_29_io_rd_data_valid; // @[pe.scala 303:15]
  wire [127:0] MemController_29_io_rd_data_bits; // @[pe.scala 303:15]
  wire  MemController_29_io_wr_data_valid; // @[pe.scala 303:15]
  wire [127:0] MemController_29_io_wr_data_bits; // @[pe.scala 303:15]
  wire  MemController_30_clock; // @[pe.scala 303:15]
  wire  MemController_30_reset; // @[pe.scala 303:15]
  wire  MemController_30_io_rd_valid; // @[pe.scala 303:15]
  wire  MemController_30_io_wr_valid; // @[pe.scala 303:15]
  wire  MemController_30_io_rd_data_valid; // @[pe.scala 303:15]
  wire [127:0] MemController_30_io_rd_data_bits; // @[pe.scala 303:15]
  wire  MemController_30_io_wr_data_valid; // @[pe.scala 303:15]
  wire [127:0] MemController_30_io_wr_data_bits; // @[pe.scala 303:15]
  wire  MemController_31_clock; // @[pe.scala 303:15]
  wire  MemController_31_reset; // @[pe.scala 303:15]
  wire  MemController_31_io_rd_valid; // @[pe.scala 303:15]
  wire  MemController_31_io_wr_valid; // @[pe.scala 303:15]
  wire  MemController_31_io_rd_data_valid; // @[pe.scala 303:15]
  wire [127:0] MemController_31_io_rd_data_bits; // @[pe.scala 303:15]
  wire  MemController_31_io_wr_data_valid; // @[pe.scala 303:15]
  wire [127:0] MemController_31_io_wr_data_bits; // @[pe.scala 303:15]
  wire  MemController_32_clock; // @[pe.scala 303:15]
  wire  MemController_32_reset; // @[pe.scala 303:15]
  wire  MemController_32_io_rd_valid; // @[pe.scala 303:15]
  wire  MemController_32_io_wr_valid; // @[pe.scala 303:15]
  wire  MemController_32_io_rd_data_valid; // @[pe.scala 303:15]
  wire [127:0] MemController_32_io_rd_data_bits; // @[pe.scala 303:15]
  wire  MemController_32_io_wr_data_valid; // @[pe.scala 303:15]
  wire [127:0] MemController_32_io_wr_data_bits; // @[pe.scala 303:15]
  wire  MemController_33_clock; // @[pe.scala 303:15]
  wire  MemController_33_reset; // @[pe.scala 303:15]
  wire  MemController_33_io_rd_valid; // @[pe.scala 303:15]
  wire  MemController_33_io_wr_valid; // @[pe.scala 303:15]
  wire  MemController_33_io_rd_data_valid; // @[pe.scala 303:15]
  wire [127:0] MemController_33_io_rd_data_bits; // @[pe.scala 303:15]
  wire  MemController_33_io_wr_data_valid; // @[pe.scala 303:15]
  wire [127:0] MemController_33_io_wr_data_bits; // @[pe.scala 303:15]
  wire  MemController_34_clock; // @[pe.scala 303:15]
  wire  MemController_34_reset; // @[pe.scala 303:15]
  wire  MemController_34_io_rd_valid; // @[pe.scala 303:15]
  wire  MemController_34_io_wr_valid; // @[pe.scala 303:15]
  wire  MemController_34_io_rd_data_valid; // @[pe.scala 303:15]
  wire [127:0] MemController_34_io_rd_data_bits; // @[pe.scala 303:15]
  wire  MemController_34_io_wr_data_valid; // @[pe.scala 303:15]
  wire [127:0] MemController_34_io_wr_data_bits; // @[pe.scala 303:15]
  wire  MemController_35_clock; // @[pe.scala 303:15]
  wire  MemController_35_reset; // @[pe.scala 303:15]
  wire  MemController_35_io_rd_valid; // @[pe.scala 303:15]
  wire  MemController_35_io_wr_valid; // @[pe.scala 303:15]
  wire  MemController_35_io_rd_data_valid; // @[pe.scala 303:15]
  wire [127:0] MemController_35_io_rd_data_bits; // @[pe.scala 303:15]
  wire  MemController_35_io_wr_data_valid; // @[pe.scala 303:15]
  wire [127:0] MemController_35_io_wr_data_bits; // @[pe.scala 303:15]
  wire  MemController_36_clock; // @[pe.scala 303:15]
  wire  MemController_36_reset; // @[pe.scala 303:15]
  wire  MemController_36_io_rd_valid; // @[pe.scala 303:15]
  wire  MemController_36_io_wr_valid; // @[pe.scala 303:15]
  wire  MemController_36_io_rd_data_valid; // @[pe.scala 303:15]
  wire [127:0] MemController_36_io_rd_data_bits; // @[pe.scala 303:15]
  wire  MemController_36_io_wr_data_valid; // @[pe.scala 303:15]
  wire [127:0] MemController_36_io_wr_data_bits; // @[pe.scala 303:15]
  wire  MemController_37_clock; // @[pe.scala 303:15]
  wire  MemController_37_reset; // @[pe.scala 303:15]
  wire  MemController_37_io_rd_valid; // @[pe.scala 303:15]
  wire  MemController_37_io_wr_valid; // @[pe.scala 303:15]
  wire  MemController_37_io_rd_data_valid; // @[pe.scala 303:15]
  wire [127:0] MemController_37_io_rd_data_bits; // @[pe.scala 303:15]
  wire  MemController_37_io_wr_data_valid; // @[pe.scala 303:15]
  wire [127:0] MemController_37_io_wr_data_bits; // @[pe.scala 303:15]
  wire  MemController_38_clock; // @[pe.scala 303:15]
  wire  MemController_38_reset; // @[pe.scala 303:15]
  wire  MemController_38_io_rd_valid; // @[pe.scala 303:15]
  wire  MemController_38_io_wr_valid; // @[pe.scala 303:15]
  wire  MemController_38_io_rd_data_valid; // @[pe.scala 303:15]
  wire [127:0] MemController_38_io_rd_data_bits; // @[pe.scala 303:15]
  wire  MemController_38_io_wr_data_valid; // @[pe.scala 303:15]
  wire [127:0] MemController_38_io_wr_data_bits; // @[pe.scala 303:15]
  wire  MemController_39_clock; // @[pe.scala 303:15]
  wire  MemController_39_reset; // @[pe.scala 303:15]
  wire  MemController_39_io_rd_valid; // @[pe.scala 303:15]
  wire  MemController_39_io_wr_valid; // @[pe.scala 303:15]
  wire  MemController_39_io_rd_data_valid; // @[pe.scala 303:15]
  wire [127:0] MemController_39_io_rd_data_bits; // @[pe.scala 303:15]
  wire  MemController_39_io_wr_data_valid; // @[pe.scala 303:15]
  wire [127:0] MemController_39_io_wr_data_bits; // @[pe.scala 303:15]
  wire  MemController_40_clock; // @[pe.scala 303:15]
  wire  MemController_40_reset; // @[pe.scala 303:15]
  wire  MemController_40_io_rd_valid; // @[pe.scala 303:15]
  wire  MemController_40_io_wr_valid; // @[pe.scala 303:15]
  wire  MemController_40_io_rd_data_valid; // @[pe.scala 303:15]
  wire [127:0] MemController_40_io_rd_data_bits; // @[pe.scala 303:15]
  wire  MemController_40_io_wr_data_valid; // @[pe.scala 303:15]
  wire [127:0] MemController_40_io_wr_data_bits; // @[pe.scala 303:15]
  wire  MemController_41_clock; // @[pe.scala 303:15]
  wire  MemController_41_reset; // @[pe.scala 303:15]
  wire  MemController_41_io_rd_valid; // @[pe.scala 303:15]
  wire  MemController_41_io_wr_valid; // @[pe.scala 303:15]
  wire  MemController_41_io_rd_data_valid; // @[pe.scala 303:15]
  wire [127:0] MemController_41_io_rd_data_bits; // @[pe.scala 303:15]
  wire  MemController_41_io_wr_data_valid; // @[pe.scala 303:15]
  wire [127:0] MemController_41_io_wr_data_bits; // @[pe.scala 303:15]
  wire  MemController_42_clock; // @[pe.scala 303:15]
  wire  MemController_42_reset; // @[pe.scala 303:15]
  wire  MemController_42_io_rd_valid; // @[pe.scala 303:15]
  wire  MemController_42_io_wr_valid; // @[pe.scala 303:15]
  wire  MemController_42_io_rd_data_valid; // @[pe.scala 303:15]
  wire [127:0] MemController_42_io_rd_data_bits; // @[pe.scala 303:15]
  wire  MemController_42_io_wr_data_valid; // @[pe.scala 303:15]
  wire [127:0] MemController_42_io_wr_data_bits; // @[pe.scala 303:15]
  wire  MemController_43_clock; // @[pe.scala 303:15]
  wire  MemController_43_reset; // @[pe.scala 303:15]
  wire  MemController_43_io_rd_valid; // @[pe.scala 303:15]
  wire  MemController_43_io_wr_valid; // @[pe.scala 303:15]
  wire  MemController_43_io_rd_data_valid; // @[pe.scala 303:15]
  wire [127:0] MemController_43_io_rd_data_bits; // @[pe.scala 303:15]
  wire  MemController_43_io_wr_data_valid; // @[pe.scala 303:15]
  wire [127:0] MemController_43_io_wr_data_bits; // @[pe.scala 303:15]
  wire  MemController_44_clock; // @[pe.scala 303:15]
  wire  MemController_44_reset; // @[pe.scala 303:15]
  wire  MemController_44_io_rd_valid; // @[pe.scala 303:15]
  wire  MemController_44_io_wr_valid; // @[pe.scala 303:15]
  wire  MemController_44_io_rd_data_valid; // @[pe.scala 303:15]
  wire [127:0] MemController_44_io_rd_data_bits; // @[pe.scala 303:15]
  wire  MemController_44_io_wr_data_valid; // @[pe.scala 303:15]
  wire [127:0] MemController_44_io_wr_data_bits; // @[pe.scala 303:15]
  wire  MemController_45_clock; // @[pe.scala 303:15]
  wire  MemController_45_reset; // @[pe.scala 303:15]
  wire  MemController_45_io_rd_valid; // @[pe.scala 303:15]
  wire  MemController_45_io_wr_valid; // @[pe.scala 303:15]
  wire  MemController_45_io_rd_data_valid; // @[pe.scala 303:15]
  wire [127:0] MemController_45_io_rd_data_bits; // @[pe.scala 303:15]
  wire  MemController_45_io_wr_data_valid; // @[pe.scala 303:15]
  wire [127:0] MemController_45_io_wr_data_bits; // @[pe.scala 303:15]
  wire  MemController_46_clock; // @[pe.scala 303:15]
  wire  MemController_46_reset; // @[pe.scala 303:15]
  wire  MemController_46_io_rd_valid; // @[pe.scala 303:15]
  wire  MemController_46_io_wr_valid; // @[pe.scala 303:15]
  wire  MemController_46_io_rd_data_valid; // @[pe.scala 303:15]
  wire [127:0] MemController_46_io_rd_data_bits; // @[pe.scala 303:15]
  wire  MemController_46_io_wr_data_valid; // @[pe.scala 303:15]
  wire [127:0] MemController_46_io_wr_data_bits; // @[pe.scala 303:15]
  wire  MemController_47_clock; // @[pe.scala 303:15]
  wire  MemController_47_reset; // @[pe.scala 303:15]
  wire  MemController_47_io_rd_valid; // @[pe.scala 303:15]
  wire  MemController_47_io_wr_valid; // @[pe.scala 303:15]
  wire  MemController_47_io_rd_data_valid; // @[pe.scala 303:15]
  wire [127:0] MemController_47_io_rd_data_bits; // @[pe.scala 303:15]
  wire  MemController_47_io_wr_data_valid; // @[pe.scala 303:15]
  wire [127:0] MemController_47_io_wr_data_bits; // @[pe.scala 303:15]
  wire  MemController_48_clock; // @[pe.scala 303:15]
  wire  MemController_48_reset; // @[pe.scala 303:15]
  wire  MemController_48_io_rd_valid; // @[pe.scala 303:15]
  wire  MemController_48_io_wr_valid; // @[pe.scala 303:15]
  wire  MemController_48_io_rd_data_valid; // @[pe.scala 303:15]
  wire [127:0] MemController_48_io_rd_data_bits; // @[pe.scala 303:15]
  wire  MemController_48_io_wr_data_valid; // @[pe.scala 303:15]
  wire [127:0] MemController_48_io_wr_data_bits; // @[pe.scala 303:15]
  wire  MemController_49_clock; // @[pe.scala 303:15]
  wire  MemController_49_reset; // @[pe.scala 303:15]
  wire  MemController_49_io_rd_valid; // @[pe.scala 303:15]
  wire  MemController_49_io_wr_valid; // @[pe.scala 303:15]
  wire  MemController_49_io_rd_data_valid; // @[pe.scala 303:15]
  wire [127:0] MemController_49_io_rd_data_bits; // @[pe.scala 303:15]
  wire  MemController_49_io_wr_data_valid; // @[pe.scala 303:15]
  wire [127:0] MemController_49_io_wr_data_bits; // @[pe.scala 303:15]
  wire  MemController_50_clock; // @[pe.scala 303:15]
  wire  MemController_50_reset; // @[pe.scala 303:15]
  wire  MemController_50_io_rd_valid; // @[pe.scala 303:15]
  wire  MemController_50_io_wr_valid; // @[pe.scala 303:15]
  wire  MemController_50_io_rd_data_valid; // @[pe.scala 303:15]
  wire [127:0] MemController_50_io_rd_data_bits; // @[pe.scala 303:15]
  wire  MemController_50_io_wr_data_valid; // @[pe.scala 303:15]
  wire [127:0] MemController_50_io_wr_data_bits; // @[pe.scala 303:15]
  wire  MemController_51_clock; // @[pe.scala 303:15]
  wire  MemController_51_reset; // @[pe.scala 303:15]
  wire  MemController_51_io_rd_valid; // @[pe.scala 303:15]
  wire  MemController_51_io_wr_valid; // @[pe.scala 303:15]
  wire  MemController_51_io_rd_data_valid; // @[pe.scala 303:15]
  wire [127:0] MemController_51_io_rd_data_bits; // @[pe.scala 303:15]
  wire  MemController_51_io_wr_data_valid; // @[pe.scala 303:15]
  wire [127:0] MemController_51_io_wr_data_bits; // @[pe.scala 303:15]
  wire  MemController_52_clock; // @[pe.scala 301:15]
  wire  MemController_52_reset; // @[pe.scala 301:15]
  wire  MemController_52_io_rd_valid; // @[pe.scala 301:15]
  wire  MemController_52_io_wr_valid; // @[pe.scala 301:15]
  wire  MemController_52_io_rd_data_valid; // @[pe.scala 301:15]
  wire [127:0] MemController_52_io_rd_data_bits; // @[pe.scala 301:15]
  wire  MemController_52_io_wr_data_valid; // @[pe.scala 301:15]
  wire [127:0] MemController_52_io_wr_data_bits; // @[pe.scala 301:15]
  wire  MemController_53_clock; // @[pe.scala 301:15]
  wire  MemController_53_reset; // @[pe.scala 301:15]
  wire  MemController_53_io_rd_valid; // @[pe.scala 301:15]
  wire  MemController_53_io_wr_valid; // @[pe.scala 301:15]
  wire  MemController_53_io_rd_data_valid; // @[pe.scala 301:15]
  wire [127:0] MemController_53_io_rd_data_bits; // @[pe.scala 301:15]
  wire  MemController_53_io_wr_data_valid; // @[pe.scala 301:15]
  wire [127:0] MemController_53_io_wr_data_bits; // @[pe.scala 301:15]
  wire  MemController_54_clock; // @[pe.scala 301:15]
  wire  MemController_54_reset; // @[pe.scala 301:15]
  wire  MemController_54_io_rd_valid; // @[pe.scala 301:15]
  wire  MemController_54_io_wr_valid; // @[pe.scala 301:15]
  wire  MemController_54_io_rd_data_valid; // @[pe.scala 301:15]
  wire [127:0] MemController_54_io_rd_data_bits; // @[pe.scala 301:15]
  wire  MemController_54_io_wr_data_valid; // @[pe.scala 301:15]
  wire [127:0] MemController_54_io_wr_data_bits; // @[pe.scala 301:15]
  wire  MemController_55_clock; // @[pe.scala 301:15]
  wire  MemController_55_reset; // @[pe.scala 301:15]
  wire  MemController_55_io_rd_valid; // @[pe.scala 301:15]
  wire  MemController_55_io_wr_valid; // @[pe.scala 301:15]
  wire  MemController_55_io_rd_data_valid; // @[pe.scala 301:15]
  wire [127:0] MemController_55_io_rd_data_bits; // @[pe.scala 301:15]
  wire  MemController_55_io_wr_data_valid; // @[pe.scala 301:15]
  wire [127:0] MemController_55_io_wr_data_bits; // @[pe.scala 301:15]
  wire  MemController_56_clock; // @[pe.scala 301:15]
  wire  MemController_56_reset; // @[pe.scala 301:15]
  wire  MemController_56_io_rd_valid; // @[pe.scala 301:15]
  wire  MemController_56_io_wr_valid; // @[pe.scala 301:15]
  wire  MemController_56_io_rd_data_valid; // @[pe.scala 301:15]
  wire [127:0] MemController_56_io_rd_data_bits; // @[pe.scala 301:15]
  wire  MemController_56_io_wr_data_valid; // @[pe.scala 301:15]
  wire [127:0] MemController_56_io_wr_data_bits; // @[pe.scala 301:15]
  wire  MemController_57_clock; // @[pe.scala 301:15]
  wire  MemController_57_reset; // @[pe.scala 301:15]
  wire  MemController_57_io_rd_valid; // @[pe.scala 301:15]
  wire  MemController_57_io_wr_valid; // @[pe.scala 301:15]
  wire  MemController_57_io_rd_data_valid; // @[pe.scala 301:15]
  wire [127:0] MemController_57_io_rd_data_bits; // @[pe.scala 301:15]
  wire  MemController_57_io_wr_data_valid; // @[pe.scala 301:15]
  wire [127:0] MemController_57_io_wr_data_bits; // @[pe.scala 301:15]
  wire  MemController_58_clock; // @[pe.scala 301:15]
  wire  MemController_58_reset; // @[pe.scala 301:15]
  wire  MemController_58_io_rd_valid; // @[pe.scala 301:15]
  wire  MemController_58_io_wr_valid; // @[pe.scala 301:15]
  wire  MemController_58_io_rd_data_valid; // @[pe.scala 301:15]
  wire [127:0] MemController_58_io_rd_data_bits; // @[pe.scala 301:15]
  wire  MemController_58_io_wr_data_valid; // @[pe.scala 301:15]
  wire [127:0] MemController_58_io_wr_data_bits; // @[pe.scala 301:15]
  wire  MemController_59_clock; // @[pe.scala 301:15]
  wire  MemController_59_reset; // @[pe.scala 301:15]
  wire  MemController_59_io_rd_valid; // @[pe.scala 301:15]
  wire  MemController_59_io_wr_valid; // @[pe.scala 301:15]
  wire  MemController_59_io_rd_data_valid; // @[pe.scala 301:15]
  wire [127:0] MemController_59_io_rd_data_bits; // @[pe.scala 301:15]
  wire  MemController_59_io_wr_data_valid; // @[pe.scala 301:15]
  wire [127:0] MemController_59_io_wr_data_bits; // @[pe.scala 301:15]
  wire  MemController_60_clock; // @[pe.scala 301:15]
  wire  MemController_60_reset; // @[pe.scala 301:15]
  wire  MemController_60_io_rd_valid; // @[pe.scala 301:15]
  wire  MemController_60_io_wr_valid; // @[pe.scala 301:15]
  wire  MemController_60_io_rd_data_valid; // @[pe.scala 301:15]
  wire [127:0] MemController_60_io_rd_data_bits; // @[pe.scala 301:15]
  wire  MemController_60_io_wr_data_valid; // @[pe.scala 301:15]
  wire [127:0] MemController_60_io_wr_data_bits; // @[pe.scala 301:15]
  wire  MemController_61_clock; // @[pe.scala 301:15]
  wire  MemController_61_reset; // @[pe.scala 301:15]
  wire  MemController_61_io_rd_valid; // @[pe.scala 301:15]
  wire  MemController_61_io_wr_valid; // @[pe.scala 301:15]
  wire  MemController_61_io_rd_data_valid; // @[pe.scala 301:15]
  wire [127:0] MemController_61_io_rd_data_bits; // @[pe.scala 301:15]
  wire  MemController_61_io_wr_data_valid; // @[pe.scala 301:15]
  wire [127:0] MemController_61_io_wr_data_bits; // @[pe.scala 301:15]
  wire  MemController_62_clock; // @[pe.scala 301:15]
  wire  MemController_62_reset; // @[pe.scala 301:15]
  wire  MemController_62_io_rd_valid; // @[pe.scala 301:15]
  wire  MemController_62_io_wr_valid; // @[pe.scala 301:15]
  wire  MemController_62_io_rd_data_valid; // @[pe.scala 301:15]
  wire [127:0] MemController_62_io_rd_data_bits; // @[pe.scala 301:15]
  wire  MemController_62_io_wr_data_valid; // @[pe.scala 301:15]
  wire [127:0] MemController_62_io_wr_data_bits; // @[pe.scala 301:15]
  wire  MemController_63_clock; // @[pe.scala 301:15]
  wire  MemController_63_reset; // @[pe.scala 301:15]
  wire  MemController_63_io_rd_valid; // @[pe.scala 301:15]
  wire  MemController_63_io_wr_valid; // @[pe.scala 301:15]
  wire  MemController_63_io_rd_data_valid; // @[pe.scala 301:15]
  wire [127:0] MemController_63_io_rd_data_bits; // @[pe.scala 301:15]
  wire  MemController_63_io_wr_data_valid; // @[pe.scala 301:15]
  wire [127:0] MemController_63_io_wr_data_bits; // @[pe.scala 301:15]
  wire  MemController_64_clock; // @[pe.scala 301:15]
  wire  MemController_64_reset; // @[pe.scala 301:15]
  wire  MemController_64_io_rd_valid; // @[pe.scala 301:15]
  wire  MemController_64_io_wr_valid; // @[pe.scala 301:15]
  wire  MemController_64_io_rd_data_valid; // @[pe.scala 301:15]
  wire [127:0] MemController_64_io_rd_data_bits; // @[pe.scala 301:15]
  wire  MemController_64_io_wr_data_valid; // @[pe.scala 301:15]
  wire [127:0] MemController_64_io_wr_data_bits; // @[pe.scala 301:15]
  wire  MemController_65_clock; // @[pe.scala 301:15]
  wire  MemController_65_reset; // @[pe.scala 301:15]
  wire  MemController_65_io_rd_valid; // @[pe.scala 301:15]
  wire  MemController_65_io_wr_valid; // @[pe.scala 301:15]
  wire  MemController_65_io_rd_data_valid; // @[pe.scala 301:15]
  wire [127:0] MemController_65_io_rd_data_bits; // @[pe.scala 301:15]
  wire  MemController_65_io_wr_data_valid; // @[pe.scala 301:15]
  wire [127:0] MemController_65_io_wr_data_bits; // @[pe.scala 301:15]
  wire  MemController_66_clock; // @[pe.scala 301:15]
  wire  MemController_66_reset; // @[pe.scala 301:15]
  wire  MemController_66_io_rd_valid; // @[pe.scala 301:15]
  wire  MemController_66_io_wr_valid; // @[pe.scala 301:15]
  wire  MemController_66_io_rd_data_valid; // @[pe.scala 301:15]
  wire [127:0] MemController_66_io_rd_data_bits; // @[pe.scala 301:15]
  wire  MemController_66_io_wr_data_valid; // @[pe.scala 301:15]
  wire [127:0] MemController_66_io_wr_data_bits; // @[pe.scala 301:15]
  wire  MemController_67_clock; // @[pe.scala 301:15]
  wire  MemController_67_reset; // @[pe.scala 301:15]
  wire  MemController_67_io_rd_valid; // @[pe.scala 301:15]
  wire  MemController_67_io_wr_valid; // @[pe.scala 301:15]
  wire  MemController_67_io_rd_data_valid; // @[pe.scala 301:15]
  wire [127:0] MemController_67_io_rd_data_bits; // @[pe.scala 301:15]
  wire  MemController_67_io_wr_data_valid; // @[pe.scala 301:15]
  wire [127:0] MemController_67_io_wr_data_bits; // @[pe.scala 301:15]
  wire  MemController_68_clock; // @[pe.scala 301:15]
  wire  MemController_68_reset; // @[pe.scala 301:15]
  wire  MemController_68_io_rd_valid; // @[pe.scala 301:15]
  wire  MemController_68_io_wr_valid; // @[pe.scala 301:15]
  wire  MemController_68_io_rd_data_valid; // @[pe.scala 301:15]
  wire [127:0] MemController_68_io_rd_data_bits; // @[pe.scala 301:15]
  wire  MemController_68_io_wr_data_valid; // @[pe.scala 301:15]
  wire [127:0] MemController_68_io_wr_data_bits; // @[pe.scala 301:15]
  wire  MemController_69_clock; // @[pe.scala 301:15]
  wire  MemController_69_reset; // @[pe.scala 301:15]
  wire  MemController_69_io_rd_valid; // @[pe.scala 301:15]
  wire  MemController_69_io_wr_valid; // @[pe.scala 301:15]
  wire  MemController_69_io_rd_data_valid; // @[pe.scala 301:15]
  wire [127:0] MemController_69_io_rd_data_bits; // @[pe.scala 301:15]
  wire  MemController_69_io_wr_data_valid; // @[pe.scala 301:15]
  wire [127:0] MemController_69_io_wr_data_bits; // @[pe.scala 301:15]
  wire  MemController_70_clock; // @[pe.scala 301:15]
  wire  MemController_70_reset; // @[pe.scala 301:15]
  wire  MemController_70_io_rd_valid; // @[pe.scala 301:15]
  wire  MemController_70_io_wr_valid; // @[pe.scala 301:15]
  wire  MemController_70_io_rd_data_valid; // @[pe.scala 301:15]
  wire [127:0] MemController_70_io_rd_data_bits; // @[pe.scala 301:15]
  wire  MemController_70_io_wr_data_valid; // @[pe.scala 301:15]
  wire [127:0] MemController_70_io_wr_data_bits; // @[pe.scala 301:15]
  wire  MemController_71_clock; // @[pe.scala 301:15]
  wire  MemController_71_reset; // @[pe.scala 301:15]
  wire  MemController_71_io_rd_valid; // @[pe.scala 301:15]
  wire  MemController_71_io_wr_valid; // @[pe.scala 301:15]
  wire  MemController_71_io_rd_data_valid; // @[pe.scala 301:15]
  wire [127:0] MemController_71_io_rd_data_bits; // @[pe.scala 301:15]
  wire  MemController_71_io_wr_data_valid; // @[pe.scala 301:15]
  wire [127:0] MemController_71_io_wr_data_bits; // @[pe.scala 301:15]
  wire  MemController_72_clock; // @[pe.scala 301:15]
  wire  MemController_72_reset; // @[pe.scala 301:15]
  wire  MemController_72_io_rd_valid; // @[pe.scala 301:15]
  wire  MemController_72_io_wr_valid; // @[pe.scala 301:15]
  wire  MemController_72_io_rd_data_valid; // @[pe.scala 301:15]
  wire [127:0] MemController_72_io_rd_data_bits; // @[pe.scala 301:15]
  wire  MemController_72_io_wr_data_valid; // @[pe.scala 301:15]
  wire [127:0] MemController_72_io_wr_data_bits; // @[pe.scala 301:15]
  wire  MemController_73_clock; // @[pe.scala 301:15]
  wire  MemController_73_reset; // @[pe.scala 301:15]
  wire  MemController_73_io_rd_valid; // @[pe.scala 301:15]
  wire  MemController_73_io_wr_valid; // @[pe.scala 301:15]
  wire  MemController_73_io_rd_data_valid; // @[pe.scala 301:15]
  wire [127:0] MemController_73_io_rd_data_bits; // @[pe.scala 301:15]
  wire  MemController_73_io_wr_data_valid; // @[pe.scala 301:15]
  wire [127:0] MemController_73_io_wr_data_bits; // @[pe.scala 301:15]
  wire  MemController_74_clock; // @[pe.scala 301:15]
  wire  MemController_74_reset; // @[pe.scala 301:15]
  wire  MemController_74_io_rd_valid; // @[pe.scala 301:15]
  wire  MemController_74_io_wr_valid; // @[pe.scala 301:15]
  wire  MemController_74_io_rd_data_valid; // @[pe.scala 301:15]
  wire [127:0] MemController_74_io_rd_data_bits; // @[pe.scala 301:15]
  wire  MemController_74_io_wr_data_valid; // @[pe.scala 301:15]
  wire [127:0] MemController_74_io_wr_data_bits; // @[pe.scala 301:15]
  wire  MemController_75_clock; // @[pe.scala 301:15]
  wire  MemController_75_reset; // @[pe.scala 301:15]
  wire  MemController_75_io_rd_valid; // @[pe.scala 301:15]
  wire  MemController_75_io_wr_valid; // @[pe.scala 301:15]
  wire  MemController_75_io_rd_data_valid; // @[pe.scala 301:15]
  wire [127:0] MemController_75_io_rd_data_bits; // @[pe.scala 301:15]
  wire  MemController_75_io_wr_data_valid; // @[pe.scala 301:15]
  wire [127:0] MemController_75_io_wr_data_bits; // @[pe.scala 301:15]
  wire  MemController_76_clock; // @[pe.scala 301:15]
  wire  MemController_76_reset; // @[pe.scala 301:15]
  wire  MemController_76_io_rd_valid; // @[pe.scala 301:15]
  wire  MemController_76_io_wr_valid; // @[pe.scala 301:15]
  wire  MemController_76_io_rd_data_valid; // @[pe.scala 301:15]
  wire [127:0] MemController_76_io_rd_data_bits; // @[pe.scala 301:15]
  wire  MemController_76_io_wr_data_valid; // @[pe.scala 301:15]
  wire [127:0] MemController_76_io_wr_data_bits; // @[pe.scala 301:15]
  wire  MemController_77_clock; // @[pe.scala 301:15]
  wire  MemController_77_reset; // @[pe.scala 301:15]
  wire  MemController_77_io_rd_valid; // @[pe.scala 301:15]
  wire  MemController_77_io_wr_valid; // @[pe.scala 301:15]
  wire  MemController_77_io_rd_data_valid; // @[pe.scala 301:15]
  wire [127:0] MemController_77_io_rd_data_bits; // @[pe.scala 301:15]
  wire  MemController_77_io_wr_data_valid; // @[pe.scala 301:15]
  wire [127:0] MemController_77_io_wr_data_bits; // @[pe.scala 301:15]
  wire  MemController_78_clock; // @[pe.scala 301:15]
  wire  MemController_78_reset; // @[pe.scala 301:15]
  wire  MemController_78_io_rd_valid; // @[pe.scala 301:15]
  wire  MemController_78_io_wr_valid; // @[pe.scala 301:15]
  wire  MemController_78_io_rd_data_valid; // @[pe.scala 301:15]
  wire [127:0] MemController_78_io_rd_data_bits; // @[pe.scala 301:15]
  wire  MemController_78_io_wr_data_valid; // @[pe.scala 301:15]
  wire [127:0] MemController_78_io_wr_data_bits; // @[pe.scala 301:15]
  wire  MemController_79_clock; // @[pe.scala 301:15]
  wire  MemController_79_reset; // @[pe.scala 301:15]
  wire  MemController_79_io_rd_valid; // @[pe.scala 301:15]
  wire  MemController_79_io_wr_valid; // @[pe.scala 301:15]
  wire  MemController_79_io_rd_data_valid; // @[pe.scala 301:15]
  wire [127:0] MemController_79_io_rd_data_bits; // @[pe.scala 301:15]
  wire  MemController_79_io_wr_data_valid; // @[pe.scala 301:15]
  wire [127:0] MemController_79_io_wr_data_bits; // @[pe.scala 301:15]
  wire  MemController_80_clock; // @[pe.scala 301:15]
  wire  MemController_80_reset; // @[pe.scala 301:15]
  wire  MemController_80_io_rd_valid; // @[pe.scala 301:15]
  wire  MemController_80_io_wr_valid; // @[pe.scala 301:15]
  wire  MemController_80_io_rd_data_valid; // @[pe.scala 301:15]
  wire [127:0] MemController_80_io_rd_data_bits; // @[pe.scala 301:15]
  wire  MemController_80_io_wr_data_valid; // @[pe.scala 301:15]
  wire [127:0] MemController_80_io_wr_data_bits; // @[pe.scala 301:15]
  wire  MemController_81_clock; // @[pe.scala 301:15]
  wire  MemController_81_reset; // @[pe.scala 301:15]
  wire  MemController_81_io_rd_valid; // @[pe.scala 301:15]
  wire  MemController_81_io_wr_valid; // @[pe.scala 301:15]
  wire  MemController_81_io_rd_data_valid; // @[pe.scala 301:15]
  wire [127:0] MemController_81_io_rd_data_bits; // @[pe.scala 301:15]
  wire  MemController_81_io_wr_data_valid; // @[pe.scala 301:15]
  wire [127:0] MemController_81_io_wr_data_bits; // @[pe.scala 301:15]
  wire  _T_1 = ~reset; // @[pe.scala 166:9]
  MultiDimTime MultiDimTime ( // @[pe.scala 165:25]
    .clock(MultiDimTime_clock),
    .reset(MultiDimTime_reset),
    .io_in(MultiDimTime_io_in),
    .io_out_0(MultiDimTime_io_out_0),
    .io_out_1(MultiDimTime_io_out_1),
    .io_out_2(MultiDimTime_io_out_2),
    .io_index_0(MultiDimTime_io_index_0),
    .io_index_1(MultiDimTime_io_index_1),
    .io_index_2(MultiDimTime_io_index_2)
  );
  PE PE ( // @[pe.scala 187:13]
    .clock(PE_clock),
    .reset(PE_reset),
    .io_data_2_out_valid(PE_io_data_2_out_valid),
    .io_data_2_out_bits(PE_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_io_data_1_in_valid),
    .io_data_1_in_bits(PE_io_data_1_in_bits),
    .io_data_1_out_valid(PE_io_data_1_out_valid),
    .io_data_1_out_bits(PE_io_data_1_out_bits),
    .io_data_0_in_valid(PE_io_data_0_in_valid),
    .io_data_0_in_bits(PE_io_data_0_in_bits),
    .io_data_0_out_valid(PE_io_data_0_out_valid),
    .io_data_0_out_bits(PE_io_data_0_out_bits)
  );
  PE PE_1 ( // @[pe.scala 187:13]
    .clock(PE_1_clock),
    .reset(PE_1_reset),
    .io_data_2_out_valid(PE_1_io_data_2_out_valid),
    .io_data_2_out_bits(PE_1_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_1_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_1_io_data_1_in_valid),
    .io_data_1_in_bits(PE_1_io_data_1_in_bits),
    .io_data_1_out_valid(PE_1_io_data_1_out_valid),
    .io_data_1_out_bits(PE_1_io_data_1_out_bits),
    .io_data_0_in_valid(PE_1_io_data_0_in_valid),
    .io_data_0_in_bits(PE_1_io_data_0_in_bits),
    .io_data_0_out_valid(PE_1_io_data_0_out_valid),
    .io_data_0_out_bits(PE_1_io_data_0_out_bits)
  );
  PE PE_2 ( // @[pe.scala 187:13]
    .clock(PE_2_clock),
    .reset(PE_2_reset),
    .io_data_2_out_valid(PE_2_io_data_2_out_valid),
    .io_data_2_out_bits(PE_2_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_2_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_2_io_data_1_in_valid),
    .io_data_1_in_bits(PE_2_io_data_1_in_bits),
    .io_data_1_out_valid(PE_2_io_data_1_out_valid),
    .io_data_1_out_bits(PE_2_io_data_1_out_bits),
    .io_data_0_in_valid(PE_2_io_data_0_in_valid),
    .io_data_0_in_bits(PE_2_io_data_0_in_bits),
    .io_data_0_out_valid(PE_2_io_data_0_out_valid),
    .io_data_0_out_bits(PE_2_io_data_0_out_bits)
  );
  PE PE_3 ( // @[pe.scala 187:13]
    .clock(PE_3_clock),
    .reset(PE_3_reset),
    .io_data_2_out_valid(PE_3_io_data_2_out_valid),
    .io_data_2_out_bits(PE_3_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_3_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_3_io_data_1_in_valid),
    .io_data_1_in_bits(PE_3_io_data_1_in_bits),
    .io_data_1_out_valid(PE_3_io_data_1_out_valid),
    .io_data_1_out_bits(PE_3_io_data_1_out_bits),
    .io_data_0_in_valid(PE_3_io_data_0_in_valid),
    .io_data_0_in_bits(PE_3_io_data_0_in_bits),
    .io_data_0_out_valid(PE_3_io_data_0_out_valid),
    .io_data_0_out_bits(PE_3_io_data_0_out_bits)
  );
  PE PE_4 ( // @[pe.scala 187:13]
    .clock(PE_4_clock),
    .reset(PE_4_reset),
    .io_data_2_out_valid(PE_4_io_data_2_out_valid),
    .io_data_2_out_bits(PE_4_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_4_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_4_io_data_1_in_valid),
    .io_data_1_in_bits(PE_4_io_data_1_in_bits),
    .io_data_1_out_valid(PE_4_io_data_1_out_valid),
    .io_data_1_out_bits(PE_4_io_data_1_out_bits),
    .io_data_0_in_valid(PE_4_io_data_0_in_valid),
    .io_data_0_in_bits(PE_4_io_data_0_in_bits),
    .io_data_0_out_valid(PE_4_io_data_0_out_valid),
    .io_data_0_out_bits(PE_4_io_data_0_out_bits)
  );
  PE PE_5 ( // @[pe.scala 187:13]
    .clock(PE_5_clock),
    .reset(PE_5_reset),
    .io_data_2_out_valid(PE_5_io_data_2_out_valid),
    .io_data_2_out_bits(PE_5_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_5_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_5_io_data_1_in_valid),
    .io_data_1_in_bits(PE_5_io_data_1_in_bits),
    .io_data_1_out_valid(PE_5_io_data_1_out_valid),
    .io_data_1_out_bits(PE_5_io_data_1_out_bits),
    .io_data_0_in_valid(PE_5_io_data_0_in_valid),
    .io_data_0_in_bits(PE_5_io_data_0_in_bits),
    .io_data_0_out_valid(PE_5_io_data_0_out_valid),
    .io_data_0_out_bits(PE_5_io_data_0_out_bits)
  );
  PE PE_6 ( // @[pe.scala 187:13]
    .clock(PE_6_clock),
    .reset(PE_6_reset),
    .io_data_2_out_valid(PE_6_io_data_2_out_valid),
    .io_data_2_out_bits(PE_6_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_6_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_6_io_data_1_in_valid),
    .io_data_1_in_bits(PE_6_io_data_1_in_bits),
    .io_data_1_out_valid(PE_6_io_data_1_out_valid),
    .io_data_1_out_bits(PE_6_io_data_1_out_bits),
    .io_data_0_in_valid(PE_6_io_data_0_in_valid),
    .io_data_0_in_bits(PE_6_io_data_0_in_bits),
    .io_data_0_out_valid(PE_6_io_data_0_out_valid),
    .io_data_0_out_bits(PE_6_io_data_0_out_bits)
  );
  PE PE_7 ( // @[pe.scala 187:13]
    .clock(PE_7_clock),
    .reset(PE_7_reset),
    .io_data_2_out_valid(PE_7_io_data_2_out_valid),
    .io_data_2_out_bits(PE_7_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_7_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_7_io_data_1_in_valid),
    .io_data_1_in_bits(PE_7_io_data_1_in_bits),
    .io_data_1_out_valid(PE_7_io_data_1_out_valid),
    .io_data_1_out_bits(PE_7_io_data_1_out_bits),
    .io_data_0_in_valid(PE_7_io_data_0_in_valid),
    .io_data_0_in_bits(PE_7_io_data_0_in_bits),
    .io_data_0_out_valid(PE_7_io_data_0_out_valid),
    .io_data_0_out_bits(PE_7_io_data_0_out_bits)
  );
  PE PE_8 ( // @[pe.scala 187:13]
    .clock(PE_8_clock),
    .reset(PE_8_reset),
    .io_data_2_out_valid(PE_8_io_data_2_out_valid),
    .io_data_2_out_bits(PE_8_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_8_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_8_io_data_1_in_valid),
    .io_data_1_in_bits(PE_8_io_data_1_in_bits),
    .io_data_1_out_valid(PE_8_io_data_1_out_valid),
    .io_data_1_out_bits(PE_8_io_data_1_out_bits),
    .io_data_0_in_valid(PE_8_io_data_0_in_valid),
    .io_data_0_in_bits(PE_8_io_data_0_in_bits),
    .io_data_0_out_valid(PE_8_io_data_0_out_valid),
    .io_data_0_out_bits(PE_8_io_data_0_out_bits)
  );
  PE PE_9 ( // @[pe.scala 187:13]
    .clock(PE_9_clock),
    .reset(PE_9_reset),
    .io_data_2_out_valid(PE_9_io_data_2_out_valid),
    .io_data_2_out_bits(PE_9_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_9_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_9_io_data_1_in_valid),
    .io_data_1_in_bits(PE_9_io_data_1_in_bits),
    .io_data_1_out_valid(PE_9_io_data_1_out_valid),
    .io_data_1_out_bits(PE_9_io_data_1_out_bits),
    .io_data_0_in_valid(PE_9_io_data_0_in_valid),
    .io_data_0_in_bits(PE_9_io_data_0_in_bits),
    .io_data_0_out_valid(PE_9_io_data_0_out_valid),
    .io_data_0_out_bits(PE_9_io_data_0_out_bits)
  );
  PE PE_10 ( // @[pe.scala 187:13]
    .clock(PE_10_clock),
    .reset(PE_10_reset),
    .io_data_2_out_valid(PE_10_io_data_2_out_valid),
    .io_data_2_out_bits(PE_10_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_10_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_10_io_data_1_in_valid),
    .io_data_1_in_bits(PE_10_io_data_1_in_bits),
    .io_data_1_out_valid(PE_10_io_data_1_out_valid),
    .io_data_1_out_bits(PE_10_io_data_1_out_bits),
    .io_data_0_in_valid(PE_10_io_data_0_in_valid),
    .io_data_0_in_bits(PE_10_io_data_0_in_bits),
    .io_data_0_out_valid(PE_10_io_data_0_out_valid),
    .io_data_0_out_bits(PE_10_io_data_0_out_bits)
  );
  PE PE_11 ( // @[pe.scala 187:13]
    .clock(PE_11_clock),
    .reset(PE_11_reset),
    .io_data_2_out_valid(PE_11_io_data_2_out_valid),
    .io_data_2_out_bits(PE_11_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_11_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_11_io_data_1_in_valid),
    .io_data_1_in_bits(PE_11_io_data_1_in_bits),
    .io_data_1_out_valid(PE_11_io_data_1_out_valid),
    .io_data_1_out_bits(PE_11_io_data_1_out_bits),
    .io_data_0_in_valid(PE_11_io_data_0_in_valid),
    .io_data_0_in_bits(PE_11_io_data_0_in_bits),
    .io_data_0_out_valid(PE_11_io_data_0_out_valid),
    .io_data_0_out_bits(PE_11_io_data_0_out_bits)
  );
  PE PE_12 ( // @[pe.scala 187:13]
    .clock(PE_12_clock),
    .reset(PE_12_reset),
    .io_data_2_out_valid(PE_12_io_data_2_out_valid),
    .io_data_2_out_bits(PE_12_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_12_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_12_io_data_1_in_valid),
    .io_data_1_in_bits(PE_12_io_data_1_in_bits),
    .io_data_1_out_valid(PE_12_io_data_1_out_valid),
    .io_data_1_out_bits(PE_12_io_data_1_out_bits),
    .io_data_0_in_valid(PE_12_io_data_0_in_valid),
    .io_data_0_in_bits(PE_12_io_data_0_in_bits),
    .io_data_0_out_valid(PE_12_io_data_0_out_valid),
    .io_data_0_out_bits(PE_12_io_data_0_out_bits)
  );
  PE PE_13 ( // @[pe.scala 187:13]
    .clock(PE_13_clock),
    .reset(PE_13_reset),
    .io_data_2_out_valid(PE_13_io_data_2_out_valid),
    .io_data_2_out_bits(PE_13_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_13_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_13_io_data_1_in_valid),
    .io_data_1_in_bits(PE_13_io_data_1_in_bits),
    .io_data_1_out_valid(PE_13_io_data_1_out_valid),
    .io_data_1_out_bits(PE_13_io_data_1_out_bits),
    .io_data_0_in_valid(PE_13_io_data_0_in_valid),
    .io_data_0_in_bits(PE_13_io_data_0_in_bits),
    .io_data_0_out_valid(PE_13_io_data_0_out_valid),
    .io_data_0_out_bits(PE_13_io_data_0_out_bits)
  );
  PE PE_14 ( // @[pe.scala 187:13]
    .clock(PE_14_clock),
    .reset(PE_14_reset),
    .io_data_2_out_valid(PE_14_io_data_2_out_valid),
    .io_data_2_out_bits(PE_14_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_14_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_14_io_data_1_in_valid),
    .io_data_1_in_bits(PE_14_io_data_1_in_bits),
    .io_data_1_out_valid(PE_14_io_data_1_out_valid),
    .io_data_1_out_bits(PE_14_io_data_1_out_bits),
    .io_data_0_in_valid(PE_14_io_data_0_in_valid),
    .io_data_0_in_bits(PE_14_io_data_0_in_bits),
    .io_data_0_out_valid(PE_14_io_data_0_out_valid),
    .io_data_0_out_bits(PE_14_io_data_0_out_bits)
  );
  PE PE_15 ( // @[pe.scala 187:13]
    .clock(PE_15_clock),
    .reset(PE_15_reset),
    .io_data_2_out_valid(PE_15_io_data_2_out_valid),
    .io_data_2_out_bits(PE_15_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_15_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_15_io_data_1_in_valid),
    .io_data_1_in_bits(PE_15_io_data_1_in_bits),
    .io_data_1_out_valid(PE_15_io_data_1_out_valid),
    .io_data_1_out_bits(PE_15_io_data_1_out_bits),
    .io_data_0_in_valid(PE_15_io_data_0_in_valid),
    .io_data_0_in_bits(PE_15_io_data_0_in_bits),
    .io_data_0_out_valid(PE_15_io_data_0_out_valid),
    .io_data_0_out_bits(PE_15_io_data_0_out_bits)
  );
  PE PE_16 ( // @[pe.scala 187:13]
    .clock(PE_16_clock),
    .reset(PE_16_reset),
    .io_data_2_out_valid(PE_16_io_data_2_out_valid),
    .io_data_2_out_bits(PE_16_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_16_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_16_io_data_1_in_valid),
    .io_data_1_in_bits(PE_16_io_data_1_in_bits),
    .io_data_1_out_valid(PE_16_io_data_1_out_valid),
    .io_data_1_out_bits(PE_16_io_data_1_out_bits),
    .io_data_0_in_valid(PE_16_io_data_0_in_valid),
    .io_data_0_in_bits(PE_16_io_data_0_in_bits),
    .io_data_0_out_valid(PE_16_io_data_0_out_valid),
    .io_data_0_out_bits(PE_16_io_data_0_out_bits)
  );
  PE PE_17 ( // @[pe.scala 187:13]
    .clock(PE_17_clock),
    .reset(PE_17_reset),
    .io_data_2_out_valid(PE_17_io_data_2_out_valid),
    .io_data_2_out_bits(PE_17_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_17_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_17_io_data_1_in_valid),
    .io_data_1_in_bits(PE_17_io_data_1_in_bits),
    .io_data_1_out_valid(PE_17_io_data_1_out_valid),
    .io_data_1_out_bits(PE_17_io_data_1_out_bits),
    .io_data_0_in_valid(PE_17_io_data_0_in_valid),
    .io_data_0_in_bits(PE_17_io_data_0_in_bits),
    .io_data_0_out_valid(PE_17_io_data_0_out_valid),
    .io_data_0_out_bits(PE_17_io_data_0_out_bits)
  );
  PE PE_18 ( // @[pe.scala 187:13]
    .clock(PE_18_clock),
    .reset(PE_18_reset),
    .io_data_2_out_valid(PE_18_io_data_2_out_valid),
    .io_data_2_out_bits(PE_18_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_18_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_18_io_data_1_in_valid),
    .io_data_1_in_bits(PE_18_io_data_1_in_bits),
    .io_data_1_out_valid(PE_18_io_data_1_out_valid),
    .io_data_1_out_bits(PE_18_io_data_1_out_bits),
    .io_data_0_in_valid(PE_18_io_data_0_in_valid),
    .io_data_0_in_bits(PE_18_io_data_0_in_bits),
    .io_data_0_out_valid(PE_18_io_data_0_out_valid),
    .io_data_0_out_bits(PE_18_io_data_0_out_bits)
  );
  PE PE_19 ( // @[pe.scala 187:13]
    .clock(PE_19_clock),
    .reset(PE_19_reset),
    .io_data_2_out_valid(PE_19_io_data_2_out_valid),
    .io_data_2_out_bits(PE_19_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_19_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_19_io_data_1_in_valid),
    .io_data_1_in_bits(PE_19_io_data_1_in_bits),
    .io_data_1_out_valid(PE_19_io_data_1_out_valid),
    .io_data_1_out_bits(PE_19_io_data_1_out_bits),
    .io_data_0_in_valid(PE_19_io_data_0_in_valid),
    .io_data_0_in_bits(PE_19_io_data_0_in_bits),
    .io_data_0_out_valid(PE_19_io_data_0_out_valid),
    .io_data_0_out_bits(PE_19_io_data_0_out_bits)
  );
  PE PE_20 ( // @[pe.scala 187:13]
    .clock(PE_20_clock),
    .reset(PE_20_reset),
    .io_data_2_out_valid(PE_20_io_data_2_out_valid),
    .io_data_2_out_bits(PE_20_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_20_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_20_io_data_1_in_valid),
    .io_data_1_in_bits(PE_20_io_data_1_in_bits),
    .io_data_1_out_valid(PE_20_io_data_1_out_valid),
    .io_data_1_out_bits(PE_20_io_data_1_out_bits),
    .io_data_0_in_valid(PE_20_io_data_0_in_valid),
    .io_data_0_in_bits(PE_20_io_data_0_in_bits),
    .io_data_0_out_valid(PE_20_io_data_0_out_valid),
    .io_data_0_out_bits(PE_20_io_data_0_out_bits)
  );
  PE PE_21 ( // @[pe.scala 187:13]
    .clock(PE_21_clock),
    .reset(PE_21_reset),
    .io_data_2_out_valid(PE_21_io_data_2_out_valid),
    .io_data_2_out_bits(PE_21_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_21_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_21_io_data_1_in_valid),
    .io_data_1_in_bits(PE_21_io_data_1_in_bits),
    .io_data_1_out_valid(PE_21_io_data_1_out_valid),
    .io_data_1_out_bits(PE_21_io_data_1_out_bits),
    .io_data_0_in_valid(PE_21_io_data_0_in_valid),
    .io_data_0_in_bits(PE_21_io_data_0_in_bits),
    .io_data_0_out_valid(PE_21_io_data_0_out_valid),
    .io_data_0_out_bits(PE_21_io_data_0_out_bits)
  );
  PE PE_22 ( // @[pe.scala 187:13]
    .clock(PE_22_clock),
    .reset(PE_22_reset),
    .io_data_2_out_valid(PE_22_io_data_2_out_valid),
    .io_data_2_out_bits(PE_22_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_22_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_22_io_data_1_in_valid),
    .io_data_1_in_bits(PE_22_io_data_1_in_bits),
    .io_data_1_out_valid(PE_22_io_data_1_out_valid),
    .io_data_1_out_bits(PE_22_io_data_1_out_bits),
    .io_data_0_in_valid(PE_22_io_data_0_in_valid),
    .io_data_0_in_bits(PE_22_io_data_0_in_bits),
    .io_data_0_out_valid(PE_22_io_data_0_out_valid),
    .io_data_0_out_bits(PE_22_io_data_0_out_bits)
  );
  PE PE_23 ( // @[pe.scala 187:13]
    .clock(PE_23_clock),
    .reset(PE_23_reset),
    .io_data_2_out_valid(PE_23_io_data_2_out_valid),
    .io_data_2_out_bits(PE_23_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_23_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_23_io_data_1_in_valid),
    .io_data_1_in_bits(PE_23_io_data_1_in_bits),
    .io_data_1_out_valid(PE_23_io_data_1_out_valid),
    .io_data_1_out_bits(PE_23_io_data_1_out_bits),
    .io_data_0_in_valid(PE_23_io_data_0_in_valid),
    .io_data_0_in_bits(PE_23_io_data_0_in_bits),
    .io_data_0_out_valid(PE_23_io_data_0_out_valid),
    .io_data_0_out_bits(PE_23_io_data_0_out_bits)
  );
  PE PE_24 ( // @[pe.scala 187:13]
    .clock(PE_24_clock),
    .reset(PE_24_reset),
    .io_data_2_out_valid(PE_24_io_data_2_out_valid),
    .io_data_2_out_bits(PE_24_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_24_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_24_io_data_1_in_valid),
    .io_data_1_in_bits(PE_24_io_data_1_in_bits),
    .io_data_1_out_valid(PE_24_io_data_1_out_valid),
    .io_data_1_out_bits(PE_24_io_data_1_out_bits),
    .io_data_0_in_valid(PE_24_io_data_0_in_valid),
    .io_data_0_in_bits(PE_24_io_data_0_in_bits),
    .io_data_0_out_valid(PE_24_io_data_0_out_valid),
    .io_data_0_out_bits(PE_24_io_data_0_out_bits)
  );
  PE PE_25 ( // @[pe.scala 187:13]
    .clock(PE_25_clock),
    .reset(PE_25_reset),
    .io_data_2_out_valid(PE_25_io_data_2_out_valid),
    .io_data_2_out_bits(PE_25_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_25_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_25_io_data_1_in_valid),
    .io_data_1_in_bits(PE_25_io_data_1_in_bits),
    .io_data_1_out_valid(PE_25_io_data_1_out_valid),
    .io_data_1_out_bits(PE_25_io_data_1_out_bits),
    .io_data_0_in_valid(PE_25_io_data_0_in_valid),
    .io_data_0_in_bits(PE_25_io_data_0_in_bits),
    .io_data_0_out_valid(PE_25_io_data_0_out_valid),
    .io_data_0_out_bits(PE_25_io_data_0_out_bits)
  );
  PE PE_26 ( // @[pe.scala 187:13]
    .clock(PE_26_clock),
    .reset(PE_26_reset),
    .io_data_2_out_valid(PE_26_io_data_2_out_valid),
    .io_data_2_out_bits(PE_26_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_26_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_26_io_data_1_in_valid),
    .io_data_1_in_bits(PE_26_io_data_1_in_bits),
    .io_data_1_out_valid(PE_26_io_data_1_out_valid),
    .io_data_1_out_bits(PE_26_io_data_1_out_bits),
    .io_data_0_in_valid(PE_26_io_data_0_in_valid),
    .io_data_0_in_bits(PE_26_io_data_0_in_bits),
    .io_data_0_out_valid(PE_26_io_data_0_out_valid),
    .io_data_0_out_bits(PE_26_io_data_0_out_bits)
  );
  PE PE_27 ( // @[pe.scala 187:13]
    .clock(PE_27_clock),
    .reset(PE_27_reset),
    .io_data_2_out_valid(PE_27_io_data_2_out_valid),
    .io_data_2_out_bits(PE_27_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_27_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_27_io_data_1_in_valid),
    .io_data_1_in_bits(PE_27_io_data_1_in_bits),
    .io_data_1_out_valid(PE_27_io_data_1_out_valid),
    .io_data_1_out_bits(PE_27_io_data_1_out_bits),
    .io_data_0_in_valid(PE_27_io_data_0_in_valid),
    .io_data_0_in_bits(PE_27_io_data_0_in_bits),
    .io_data_0_out_valid(PE_27_io_data_0_out_valid),
    .io_data_0_out_bits(PE_27_io_data_0_out_bits)
  );
  PE PE_28 ( // @[pe.scala 187:13]
    .clock(PE_28_clock),
    .reset(PE_28_reset),
    .io_data_2_out_valid(PE_28_io_data_2_out_valid),
    .io_data_2_out_bits(PE_28_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_28_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_28_io_data_1_in_valid),
    .io_data_1_in_bits(PE_28_io_data_1_in_bits),
    .io_data_1_out_valid(PE_28_io_data_1_out_valid),
    .io_data_1_out_bits(PE_28_io_data_1_out_bits),
    .io_data_0_in_valid(PE_28_io_data_0_in_valid),
    .io_data_0_in_bits(PE_28_io_data_0_in_bits),
    .io_data_0_out_valid(PE_28_io_data_0_out_valid),
    .io_data_0_out_bits(PE_28_io_data_0_out_bits)
  );
  PE PE_29 ( // @[pe.scala 187:13]
    .clock(PE_29_clock),
    .reset(PE_29_reset),
    .io_data_2_out_valid(PE_29_io_data_2_out_valid),
    .io_data_2_out_bits(PE_29_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_29_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_29_io_data_1_in_valid),
    .io_data_1_in_bits(PE_29_io_data_1_in_bits),
    .io_data_1_out_valid(PE_29_io_data_1_out_valid),
    .io_data_1_out_bits(PE_29_io_data_1_out_bits),
    .io_data_0_in_valid(PE_29_io_data_0_in_valid),
    .io_data_0_in_bits(PE_29_io_data_0_in_bits),
    .io_data_0_out_valid(PE_29_io_data_0_out_valid),
    .io_data_0_out_bits(PE_29_io_data_0_out_bits)
  );
  PE PE_30 ( // @[pe.scala 187:13]
    .clock(PE_30_clock),
    .reset(PE_30_reset),
    .io_data_2_out_valid(PE_30_io_data_2_out_valid),
    .io_data_2_out_bits(PE_30_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_30_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_30_io_data_1_in_valid),
    .io_data_1_in_bits(PE_30_io_data_1_in_bits),
    .io_data_1_out_valid(PE_30_io_data_1_out_valid),
    .io_data_1_out_bits(PE_30_io_data_1_out_bits),
    .io_data_0_in_valid(PE_30_io_data_0_in_valid),
    .io_data_0_in_bits(PE_30_io_data_0_in_bits),
    .io_data_0_out_valid(PE_30_io_data_0_out_valid),
    .io_data_0_out_bits(PE_30_io_data_0_out_bits)
  );
  PE PE_31 ( // @[pe.scala 187:13]
    .clock(PE_31_clock),
    .reset(PE_31_reset),
    .io_data_2_out_valid(PE_31_io_data_2_out_valid),
    .io_data_2_out_bits(PE_31_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_31_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_31_io_data_1_in_valid),
    .io_data_1_in_bits(PE_31_io_data_1_in_bits),
    .io_data_1_out_valid(PE_31_io_data_1_out_valid),
    .io_data_1_out_bits(PE_31_io_data_1_out_bits),
    .io_data_0_in_valid(PE_31_io_data_0_in_valid),
    .io_data_0_in_bits(PE_31_io_data_0_in_bits),
    .io_data_0_out_valid(PE_31_io_data_0_out_valid),
    .io_data_0_out_bits(PE_31_io_data_0_out_bits)
  );
  PE PE_32 ( // @[pe.scala 187:13]
    .clock(PE_32_clock),
    .reset(PE_32_reset),
    .io_data_2_out_valid(PE_32_io_data_2_out_valid),
    .io_data_2_out_bits(PE_32_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_32_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_32_io_data_1_in_valid),
    .io_data_1_in_bits(PE_32_io_data_1_in_bits),
    .io_data_1_out_valid(PE_32_io_data_1_out_valid),
    .io_data_1_out_bits(PE_32_io_data_1_out_bits),
    .io_data_0_in_valid(PE_32_io_data_0_in_valid),
    .io_data_0_in_bits(PE_32_io_data_0_in_bits),
    .io_data_0_out_valid(PE_32_io_data_0_out_valid),
    .io_data_0_out_bits(PE_32_io_data_0_out_bits)
  );
  PE PE_33 ( // @[pe.scala 187:13]
    .clock(PE_33_clock),
    .reset(PE_33_reset),
    .io_data_2_out_valid(PE_33_io_data_2_out_valid),
    .io_data_2_out_bits(PE_33_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_33_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_33_io_data_1_in_valid),
    .io_data_1_in_bits(PE_33_io_data_1_in_bits),
    .io_data_1_out_valid(PE_33_io_data_1_out_valid),
    .io_data_1_out_bits(PE_33_io_data_1_out_bits),
    .io_data_0_in_valid(PE_33_io_data_0_in_valid),
    .io_data_0_in_bits(PE_33_io_data_0_in_bits),
    .io_data_0_out_valid(PE_33_io_data_0_out_valid),
    .io_data_0_out_bits(PE_33_io_data_0_out_bits)
  );
  PE PE_34 ( // @[pe.scala 187:13]
    .clock(PE_34_clock),
    .reset(PE_34_reset),
    .io_data_2_out_valid(PE_34_io_data_2_out_valid),
    .io_data_2_out_bits(PE_34_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_34_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_34_io_data_1_in_valid),
    .io_data_1_in_bits(PE_34_io_data_1_in_bits),
    .io_data_1_out_valid(PE_34_io_data_1_out_valid),
    .io_data_1_out_bits(PE_34_io_data_1_out_bits),
    .io_data_0_in_valid(PE_34_io_data_0_in_valid),
    .io_data_0_in_bits(PE_34_io_data_0_in_bits),
    .io_data_0_out_valid(PE_34_io_data_0_out_valid),
    .io_data_0_out_bits(PE_34_io_data_0_out_bits)
  );
  PE PE_35 ( // @[pe.scala 187:13]
    .clock(PE_35_clock),
    .reset(PE_35_reset),
    .io_data_2_out_valid(PE_35_io_data_2_out_valid),
    .io_data_2_out_bits(PE_35_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_35_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_35_io_data_1_in_valid),
    .io_data_1_in_bits(PE_35_io_data_1_in_bits),
    .io_data_1_out_valid(PE_35_io_data_1_out_valid),
    .io_data_1_out_bits(PE_35_io_data_1_out_bits),
    .io_data_0_in_valid(PE_35_io_data_0_in_valid),
    .io_data_0_in_bits(PE_35_io_data_0_in_bits),
    .io_data_0_out_valid(PE_35_io_data_0_out_valid),
    .io_data_0_out_bits(PE_35_io_data_0_out_bits)
  );
  PE PE_36 ( // @[pe.scala 187:13]
    .clock(PE_36_clock),
    .reset(PE_36_reset),
    .io_data_2_out_valid(PE_36_io_data_2_out_valid),
    .io_data_2_out_bits(PE_36_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_36_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_36_io_data_1_in_valid),
    .io_data_1_in_bits(PE_36_io_data_1_in_bits),
    .io_data_1_out_valid(PE_36_io_data_1_out_valid),
    .io_data_1_out_bits(PE_36_io_data_1_out_bits),
    .io_data_0_in_valid(PE_36_io_data_0_in_valid),
    .io_data_0_in_bits(PE_36_io_data_0_in_bits),
    .io_data_0_out_valid(PE_36_io_data_0_out_valid),
    .io_data_0_out_bits(PE_36_io_data_0_out_bits)
  );
  PE PE_37 ( // @[pe.scala 187:13]
    .clock(PE_37_clock),
    .reset(PE_37_reset),
    .io_data_2_out_valid(PE_37_io_data_2_out_valid),
    .io_data_2_out_bits(PE_37_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_37_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_37_io_data_1_in_valid),
    .io_data_1_in_bits(PE_37_io_data_1_in_bits),
    .io_data_1_out_valid(PE_37_io_data_1_out_valid),
    .io_data_1_out_bits(PE_37_io_data_1_out_bits),
    .io_data_0_in_valid(PE_37_io_data_0_in_valid),
    .io_data_0_in_bits(PE_37_io_data_0_in_bits),
    .io_data_0_out_valid(PE_37_io_data_0_out_valid),
    .io_data_0_out_bits(PE_37_io_data_0_out_bits)
  );
  PE PE_38 ( // @[pe.scala 187:13]
    .clock(PE_38_clock),
    .reset(PE_38_reset),
    .io_data_2_out_valid(PE_38_io_data_2_out_valid),
    .io_data_2_out_bits(PE_38_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_38_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_38_io_data_1_in_valid),
    .io_data_1_in_bits(PE_38_io_data_1_in_bits),
    .io_data_1_out_valid(PE_38_io_data_1_out_valid),
    .io_data_1_out_bits(PE_38_io_data_1_out_bits),
    .io_data_0_in_valid(PE_38_io_data_0_in_valid),
    .io_data_0_in_bits(PE_38_io_data_0_in_bits),
    .io_data_0_out_valid(PE_38_io_data_0_out_valid),
    .io_data_0_out_bits(PE_38_io_data_0_out_bits)
  );
  PE PE_39 ( // @[pe.scala 187:13]
    .clock(PE_39_clock),
    .reset(PE_39_reset),
    .io_data_2_out_valid(PE_39_io_data_2_out_valid),
    .io_data_2_out_bits(PE_39_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_39_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_39_io_data_1_in_valid),
    .io_data_1_in_bits(PE_39_io_data_1_in_bits),
    .io_data_1_out_valid(PE_39_io_data_1_out_valid),
    .io_data_1_out_bits(PE_39_io_data_1_out_bits),
    .io_data_0_in_valid(PE_39_io_data_0_in_valid),
    .io_data_0_in_bits(PE_39_io_data_0_in_bits),
    .io_data_0_out_valid(PE_39_io_data_0_out_valid),
    .io_data_0_out_bits(PE_39_io_data_0_out_bits)
  );
  PE PE_40 ( // @[pe.scala 187:13]
    .clock(PE_40_clock),
    .reset(PE_40_reset),
    .io_data_2_out_valid(PE_40_io_data_2_out_valid),
    .io_data_2_out_bits(PE_40_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_40_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_40_io_data_1_in_valid),
    .io_data_1_in_bits(PE_40_io_data_1_in_bits),
    .io_data_1_out_valid(PE_40_io_data_1_out_valid),
    .io_data_1_out_bits(PE_40_io_data_1_out_bits),
    .io_data_0_in_valid(PE_40_io_data_0_in_valid),
    .io_data_0_in_bits(PE_40_io_data_0_in_bits),
    .io_data_0_out_valid(PE_40_io_data_0_out_valid),
    .io_data_0_out_bits(PE_40_io_data_0_out_bits)
  );
  PE PE_41 ( // @[pe.scala 187:13]
    .clock(PE_41_clock),
    .reset(PE_41_reset),
    .io_data_2_out_valid(PE_41_io_data_2_out_valid),
    .io_data_2_out_bits(PE_41_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_41_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_41_io_data_1_in_valid),
    .io_data_1_in_bits(PE_41_io_data_1_in_bits),
    .io_data_1_out_valid(PE_41_io_data_1_out_valid),
    .io_data_1_out_bits(PE_41_io_data_1_out_bits),
    .io_data_0_in_valid(PE_41_io_data_0_in_valid),
    .io_data_0_in_bits(PE_41_io_data_0_in_bits),
    .io_data_0_out_valid(PE_41_io_data_0_out_valid),
    .io_data_0_out_bits(PE_41_io_data_0_out_bits)
  );
  PE PE_42 ( // @[pe.scala 187:13]
    .clock(PE_42_clock),
    .reset(PE_42_reset),
    .io_data_2_out_valid(PE_42_io_data_2_out_valid),
    .io_data_2_out_bits(PE_42_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_42_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_42_io_data_1_in_valid),
    .io_data_1_in_bits(PE_42_io_data_1_in_bits),
    .io_data_1_out_valid(PE_42_io_data_1_out_valid),
    .io_data_1_out_bits(PE_42_io_data_1_out_bits),
    .io_data_0_in_valid(PE_42_io_data_0_in_valid),
    .io_data_0_in_bits(PE_42_io_data_0_in_bits),
    .io_data_0_out_valid(PE_42_io_data_0_out_valid),
    .io_data_0_out_bits(PE_42_io_data_0_out_bits)
  );
  PE PE_43 ( // @[pe.scala 187:13]
    .clock(PE_43_clock),
    .reset(PE_43_reset),
    .io_data_2_out_valid(PE_43_io_data_2_out_valid),
    .io_data_2_out_bits(PE_43_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_43_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_43_io_data_1_in_valid),
    .io_data_1_in_bits(PE_43_io_data_1_in_bits),
    .io_data_1_out_valid(PE_43_io_data_1_out_valid),
    .io_data_1_out_bits(PE_43_io_data_1_out_bits),
    .io_data_0_in_valid(PE_43_io_data_0_in_valid),
    .io_data_0_in_bits(PE_43_io_data_0_in_bits),
    .io_data_0_out_valid(PE_43_io_data_0_out_valid),
    .io_data_0_out_bits(PE_43_io_data_0_out_bits)
  );
  PE PE_44 ( // @[pe.scala 187:13]
    .clock(PE_44_clock),
    .reset(PE_44_reset),
    .io_data_2_out_valid(PE_44_io_data_2_out_valid),
    .io_data_2_out_bits(PE_44_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_44_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_44_io_data_1_in_valid),
    .io_data_1_in_bits(PE_44_io_data_1_in_bits),
    .io_data_1_out_valid(PE_44_io_data_1_out_valid),
    .io_data_1_out_bits(PE_44_io_data_1_out_bits),
    .io_data_0_in_valid(PE_44_io_data_0_in_valid),
    .io_data_0_in_bits(PE_44_io_data_0_in_bits),
    .io_data_0_out_valid(PE_44_io_data_0_out_valid),
    .io_data_0_out_bits(PE_44_io_data_0_out_bits)
  );
  PE PE_45 ( // @[pe.scala 187:13]
    .clock(PE_45_clock),
    .reset(PE_45_reset),
    .io_data_2_out_valid(PE_45_io_data_2_out_valid),
    .io_data_2_out_bits(PE_45_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_45_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_45_io_data_1_in_valid),
    .io_data_1_in_bits(PE_45_io_data_1_in_bits),
    .io_data_1_out_valid(PE_45_io_data_1_out_valid),
    .io_data_1_out_bits(PE_45_io_data_1_out_bits),
    .io_data_0_in_valid(PE_45_io_data_0_in_valid),
    .io_data_0_in_bits(PE_45_io_data_0_in_bits),
    .io_data_0_out_valid(PE_45_io_data_0_out_valid),
    .io_data_0_out_bits(PE_45_io_data_0_out_bits)
  );
  PE PE_46 ( // @[pe.scala 187:13]
    .clock(PE_46_clock),
    .reset(PE_46_reset),
    .io_data_2_out_valid(PE_46_io_data_2_out_valid),
    .io_data_2_out_bits(PE_46_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_46_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_46_io_data_1_in_valid),
    .io_data_1_in_bits(PE_46_io_data_1_in_bits),
    .io_data_1_out_valid(PE_46_io_data_1_out_valid),
    .io_data_1_out_bits(PE_46_io_data_1_out_bits),
    .io_data_0_in_valid(PE_46_io_data_0_in_valid),
    .io_data_0_in_bits(PE_46_io_data_0_in_bits),
    .io_data_0_out_valid(PE_46_io_data_0_out_valid),
    .io_data_0_out_bits(PE_46_io_data_0_out_bits)
  );
  PE PE_47 ( // @[pe.scala 187:13]
    .clock(PE_47_clock),
    .reset(PE_47_reset),
    .io_data_2_out_valid(PE_47_io_data_2_out_valid),
    .io_data_2_out_bits(PE_47_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_47_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_47_io_data_1_in_valid),
    .io_data_1_in_bits(PE_47_io_data_1_in_bits),
    .io_data_1_out_valid(PE_47_io_data_1_out_valid),
    .io_data_1_out_bits(PE_47_io_data_1_out_bits),
    .io_data_0_in_valid(PE_47_io_data_0_in_valid),
    .io_data_0_in_bits(PE_47_io_data_0_in_bits),
    .io_data_0_out_valid(PE_47_io_data_0_out_valid),
    .io_data_0_out_bits(PE_47_io_data_0_out_bits)
  );
  PE PE_48 ( // @[pe.scala 187:13]
    .clock(PE_48_clock),
    .reset(PE_48_reset),
    .io_data_2_out_valid(PE_48_io_data_2_out_valid),
    .io_data_2_out_bits(PE_48_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_48_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_48_io_data_1_in_valid),
    .io_data_1_in_bits(PE_48_io_data_1_in_bits),
    .io_data_1_out_valid(PE_48_io_data_1_out_valid),
    .io_data_1_out_bits(PE_48_io_data_1_out_bits),
    .io_data_0_in_valid(PE_48_io_data_0_in_valid),
    .io_data_0_in_bits(PE_48_io_data_0_in_bits),
    .io_data_0_out_valid(PE_48_io_data_0_out_valid),
    .io_data_0_out_bits(PE_48_io_data_0_out_bits)
  );
  PE PE_49 ( // @[pe.scala 187:13]
    .clock(PE_49_clock),
    .reset(PE_49_reset),
    .io_data_2_out_valid(PE_49_io_data_2_out_valid),
    .io_data_2_out_bits(PE_49_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_49_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_49_io_data_1_in_valid),
    .io_data_1_in_bits(PE_49_io_data_1_in_bits),
    .io_data_1_out_valid(PE_49_io_data_1_out_valid),
    .io_data_1_out_bits(PE_49_io_data_1_out_bits),
    .io_data_0_in_valid(PE_49_io_data_0_in_valid),
    .io_data_0_in_bits(PE_49_io_data_0_in_bits),
    .io_data_0_out_valid(PE_49_io_data_0_out_valid),
    .io_data_0_out_bits(PE_49_io_data_0_out_bits)
  );
  PE PE_50 ( // @[pe.scala 187:13]
    .clock(PE_50_clock),
    .reset(PE_50_reset),
    .io_data_2_out_valid(PE_50_io_data_2_out_valid),
    .io_data_2_out_bits(PE_50_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_50_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_50_io_data_1_in_valid),
    .io_data_1_in_bits(PE_50_io_data_1_in_bits),
    .io_data_1_out_valid(PE_50_io_data_1_out_valid),
    .io_data_1_out_bits(PE_50_io_data_1_out_bits),
    .io_data_0_in_valid(PE_50_io_data_0_in_valid),
    .io_data_0_in_bits(PE_50_io_data_0_in_bits),
    .io_data_0_out_valid(PE_50_io_data_0_out_valid),
    .io_data_0_out_bits(PE_50_io_data_0_out_bits)
  );
  PE PE_51 ( // @[pe.scala 187:13]
    .clock(PE_51_clock),
    .reset(PE_51_reset),
    .io_data_2_out_valid(PE_51_io_data_2_out_valid),
    .io_data_2_out_bits(PE_51_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_51_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_51_io_data_1_in_valid),
    .io_data_1_in_bits(PE_51_io_data_1_in_bits),
    .io_data_1_out_valid(PE_51_io_data_1_out_valid),
    .io_data_1_out_bits(PE_51_io_data_1_out_bits),
    .io_data_0_in_valid(PE_51_io_data_0_in_valid),
    .io_data_0_in_bits(PE_51_io_data_0_in_bits),
    .io_data_0_out_valid(PE_51_io_data_0_out_valid),
    .io_data_0_out_bits(PE_51_io_data_0_out_bits)
  );
  PE PE_52 ( // @[pe.scala 187:13]
    .clock(PE_52_clock),
    .reset(PE_52_reset),
    .io_data_2_out_valid(PE_52_io_data_2_out_valid),
    .io_data_2_out_bits(PE_52_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_52_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_52_io_data_1_in_valid),
    .io_data_1_in_bits(PE_52_io_data_1_in_bits),
    .io_data_1_out_valid(PE_52_io_data_1_out_valid),
    .io_data_1_out_bits(PE_52_io_data_1_out_bits),
    .io_data_0_in_valid(PE_52_io_data_0_in_valid),
    .io_data_0_in_bits(PE_52_io_data_0_in_bits),
    .io_data_0_out_valid(PE_52_io_data_0_out_valid),
    .io_data_0_out_bits(PE_52_io_data_0_out_bits)
  );
  PE PE_53 ( // @[pe.scala 187:13]
    .clock(PE_53_clock),
    .reset(PE_53_reset),
    .io_data_2_out_valid(PE_53_io_data_2_out_valid),
    .io_data_2_out_bits(PE_53_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_53_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_53_io_data_1_in_valid),
    .io_data_1_in_bits(PE_53_io_data_1_in_bits),
    .io_data_1_out_valid(PE_53_io_data_1_out_valid),
    .io_data_1_out_bits(PE_53_io_data_1_out_bits),
    .io_data_0_in_valid(PE_53_io_data_0_in_valid),
    .io_data_0_in_bits(PE_53_io_data_0_in_bits),
    .io_data_0_out_valid(PE_53_io_data_0_out_valid),
    .io_data_0_out_bits(PE_53_io_data_0_out_bits)
  );
  PE PE_54 ( // @[pe.scala 187:13]
    .clock(PE_54_clock),
    .reset(PE_54_reset),
    .io_data_2_out_valid(PE_54_io_data_2_out_valid),
    .io_data_2_out_bits(PE_54_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_54_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_54_io_data_1_in_valid),
    .io_data_1_in_bits(PE_54_io_data_1_in_bits),
    .io_data_1_out_valid(PE_54_io_data_1_out_valid),
    .io_data_1_out_bits(PE_54_io_data_1_out_bits),
    .io_data_0_in_valid(PE_54_io_data_0_in_valid),
    .io_data_0_in_bits(PE_54_io_data_0_in_bits),
    .io_data_0_out_valid(PE_54_io_data_0_out_valid),
    .io_data_0_out_bits(PE_54_io_data_0_out_bits)
  );
  PE PE_55 ( // @[pe.scala 187:13]
    .clock(PE_55_clock),
    .reset(PE_55_reset),
    .io_data_2_out_valid(PE_55_io_data_2_out_valid),
    .io_data_2_out_bits(PE_55_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_55_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_55_io_data_1_in_valid),
    .io_data_1_in_bits(PE_55_io_data_1_in_bits),
    .io_data_1_out_valid(PE_55_io_data_1_out_valid),
    .io_data_1_out_bits(PE_55_io_data_1_out_bits),
    .io_data_0_in_valid(PE_55_io_data_0_in_valid),
    .io_data_0_in_bits(PE_55_io_data_0_in_bits),
    .io_data_0_out_valid(PE_55_io_data_0_out_valid),
    .io_data_0_out_bits(PE_55_io_data_0_out_bits)
  );
  PE PE_56 ( // @[pe.scala 187:13]
    .clock(PE_56_clock),
    .reset(PE_56_reset),
    .io_data_2_out_valid(PE_56_io_data_2_out_valid),
    .io_data_2_out_bits(PE_56_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_56_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_56_io_data_1_in_valid),
    .io_data_1_in_bits(PE_56_io_data_1_in_bits),
    .io_data_1_out_valid(PE_56_io_data_1_out_valid),
    .io_data_1_out_bits(PE_56_io_data_1_out_bits),
    .io_data_0_in_valid(PE_56_io_data_0_in_valid),
    .io_data_0_in_bits(PE_56_io_data_0_in_bits),
    .io_data_0_out_valid(PE_56_io_data_0_out_valid),
    .io_data_0_out_bits(PE_56_io_data_0_out_bits)
  );
  PE PE_57 ( // @[pe.scala 187:13]
    .clock(PE_57_clock),
    .reset(PE_57_reset),
    .io_data_2_out_valid(PE_57_io_data_2_out_valid),
    .io_data_2_out_bits(PE_57_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_57_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_57_io_data_1_in_valid),
    .io_data_1_in_bits(PE_57_io_data_1_in_bits),
    .io_data_1_out_valid(PE_57_io_data_1_out_valid),
    .io_data_1_out_bits(PE_57_io_data_1_out_bits),
    .io_data_0_in_valid(PE_57_io_data_0_in_valid),
    .io_data_0_in_bits(PE_57_io_data_0_in_bits),
    .io_data_0_out_valid(PE_57_io_data_0_out_valid),
    .io_data_0_out_bits(PE_57_io_data_0_out_bits)
  );
  PE PE_58 ( // @[pe.scala 187:13]
    .clock(PE_58_clock),
    .reset(PE_58_reset),
    .io_data_2_out_valid(PE_58_io_data_2_out_valid),
    .io_data_2_out_bits(PE_58_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_58_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_58_io_data_1_in_valid),
    .io_data_1_in_bits(PE_58_io_data_1_in_bits),
    .io_data_1_out_valid(PE_58_io_data_1_out_valid),
    .io_data_1_out_bits(PE_58_io_data_1_out_bits),
    .io_data_0_in_valid(PE_58_io_data_0_in_valid),
    .io_data_0_in_bits(PE_58_io_data_0_in_bits),
    .io_data_0_out_valid(PE_58_io_data_0_out_valid),
    .io_data_0_out_bits(PE_58_io_data_0_out_bits)
  );
  PE PE_59 ( // @[pe.scala 187:13]
    .clock(PE_59_clock),
    .reset(PE_59_reset),
    .io_data_2_out_valid(PE_59_io_data_2_out_valid),
    .io_data_2_out_bits(PE_59_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_59_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_59_io_data_1_in_valid),
    .io_data_1_in_bits(PE_59_io_data_1_in_bits),
    .io_data_1_out_valid(PE_59_io_data_1_out_valid),
    .io_data_1_out_bits(PE_59_io_data_1_out_bits),
    .io_data_0_in_valid(PE_59_io_data_0_in_valid),
    .io_data_0_in_bits(PE_59_io_data_0_in_bits),
    .io_data_0_out_valid(PE_59_io_data_0_out_valid),
    .io_data_0_out_bits(PE_59_io_data_0_out_bits)
  );
  PE PE_60 ( // @[pe.scala 187:13]
    .clock(PE_60_clock),
    .reset(PE_60_reset),
    .io_data_2_out_valid(PE_60_io_data_2_out_valid),
    .io_data_2_out_bits(PE_60_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_60_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_60_io_data_1_in_valid),
    .io_data_1_in_bits(PE_60_io_data_1_in_bits),
    .io_data_1_out_valid(PE_60_io_data_1_out_valid),
    .io_data_1_out_bits(PE_60_io_data_1_out_bits),
    .io_data_0_in_valid(PE_60_io_data_0_in_valid),
    .io_data_0_in_bits(PE_60_io_data_0_in_bits),
    .io_data_0_out_valid(PE_60_io_data_0_out_valid),
    .io_data_0_out_bits(PE_60_io_data_0_out_bits)
  );
  PE PE_61 ( // @[pe.scala 187:13]
    .clock(PE_61_clock),
    .reset(PE_61_reset),
    .io_data_2_out_valid(PE_61_io_data_2_out_valid),
    .io_data_2_out_bits(PE_61_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_61_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_61_io_data_1_in_valid),
    .io_data_1_in_bits(PE_61_io_data_1_in_bits),
    .io_data_1_out_valid(PE_61_io_data_1_out_valid),
    .io_data_1_out_bits(PE_61_io_data_1_out_bits),
    .io_data_0_in_valid(PE_61_io_data_0_in_valid),
    .io_data_0_in_bits(PE_61_io_data_0_in_bits),
    .io_data_0_out_valid(PE_61_io_data_0_out_valid),
    .io_data_0_out_bits(PE_61_io_data_0_out_bits)
  );
  PE PE_62 ( // @[pe.scala 187:13]
    .clock(PE_62_clock),
    .reset(PE_62_reset),
    .io_data_2_out_valid(PE_62_io_data_2_out_valid),
    .io_data_2_out_bits(PE_62_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_62_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_62_io_data_1_in_valid),
    .io_data_1_in_bits(PE_62_io_data_1_in_bits),
    .io_data_1_out_valid(PE_62_io_data_1_out_valid),
    .io_data_1_out_bits(PE_62_io_data_1_out_bits),
    .io_data_0_in_valid(PE_62_io_data_0_in_valid),
    .io_data_0_in_bits(PE_62_io_data_0_in_bits),
    .io_data_0_out_valid(PE_62_io_data_0_out_valid),
    .io_data_0_out_bits(PE_62_io_data_0_out_bits)
  );
  PE PE_63 ( // @[pe.scala 187:13]
    .clock(PE_63_clock),
    .reset(PE_63_reset),
    .io_data_2_out_valid(PE_63_io_data_2_out_valid),
    .io_data_2_out_bits(PE_63_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_63_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_63_io_data_1_in_valid),
    .io_data_1_in_bits(PE_63_io_data_1_in_bits),
    .io_data_1_out_valid(PE_63_io_data_1_out_valid),
    .io_data_1_out_bits(PE_63_io_data_1_out_bits),
    .io_data_0_in_valid(PE_63_io_data_0_in_valid),
    .io_data_0_in_bits(PE_63_io_data_0_in_bits),
    .io_data_0_out_valid(PE_63_io_data_0_out_valid),
    .io_data_0_out_bits(PE_63_io_data_0_out_bits)
  );
  PE PE_64 ( // @[pe.scala 187:13]
    .clock(PE_64_clock),
    .reset(PE_64_reset),
    .io_data_2_out_valid(PE_64_io_data_2_out_valid),
    .io_data_2_out_bits(PE_64_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_64_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_64_io_data_1_in_valid),
    .io_data_1_in_bits(PE_64_io_data_1_in_bits),
    .io_data_1_out_valid(PE_64_io_data_1_out_valid),
    .io_data_1_out_bits(PE_64_io_data_1_out_bits),
    .io_data_0_in_valid(PE_64_io_data_0_in_valid),
    .io_data_0_in_bits(PE_64_io_data_0_in_bits),
    .io_data_0_out_valid(PE_64_io_data_0_out_valid),
    .io_data_0_out_bits(PE_64_io_data_0_out_bits)
  );
  PE PE_65 ( // @[pe.scala 187:13]
    .clock(PE_65_clock),
    .reset(PE_65_reset),
    .io_data_2_out_valid(PE_65_io_data_2_out_valid),
    .io_data_2_out_bits(PE_65_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_65_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_65_io_data_1_in_valid),
    .io_data_1_in_bits(PE_65_io_data_1_in_bits),
    .io_data_1_out_valid(PE_65_io_data_1_out_valid),
    .io_data_1_out_bits(PE_65_io_data_1_out_bits),
    .io_data_0_in_valid(PE_65_io_data_0_in_valid),
    .io_data_0_in_bits(PE_65_io_data_0_in_bits),
    .io_data_0_out_valid(PE_65_io_data_0_out_valid),
    .io_data_0_out_bits(PE_65_io_data_0_out_bits)
  );
  PE PE_66 ( // @[pe.scala 187:13]
    .clock(PE_66_clock),
    .reset(PE_66_reset),
    .io_data_2_out_valid(PE_66_io_data_2_out_valid),
    .io_data_2_out_bits(PE_66_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_66_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_66_io_data_1_in_valid),
    .io_data_1_in_bits(PE_66_io_data_1_in_bits),
    .io_data_1_out_valid(PE_66_io_data_1_out_valid),
    .io_data_1_out_bits(PE_66_io_data_1_out_bits),
    .io_data_0_in_valid(PE_66_io_data_0_in_valid),
    .io_data_0_in_bits(PE_66_io_data_0_in_bits),
    .io_data_0_out_valid(PE_66_io_data_0_out_valid),
    .io_data_0_out_bits(PE_66_io_data_0_out_bits)
  );
  PE PE_67 ( // @[pe.scala 187:13]
    .clock(PE_67_clock),
    .reset(PE_67_reset),
    .io_data_2_out_valid(PE_67_io_data_2_out_valid),
    .io_data_2_out_bits(PE_67_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_67_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_67_io_data_1_in_valid),
    .io_data_1_in_bits(PE_67_io_data_1_in_bits),
    .io_data_1_out_valid(PE_67_io_data_1_out_valid),
    .io_data_1_out_bits(PE_67_io_data_1_out_bits),
    .io_data_0_in_valid(PE_67_io_data_0_in_valid),
    .io_data_0_in_bits(PE_67_io_data_0_in_bits),
    .io_data_0_out_valid(PE_67_io_data_0_out_valid),
    .io_data_0_out_bits(PE_67_io_data_0_out_bits)
  );
  PE PE_68 ( // @[pe.scala 187:13]
    .clock(PE_68_clock),
    .reset(PE_68_reset),
    .io_data_2_out_valid(PE_68_io_data_2_out_valid),
    .io_data_2_out_bits(PE_68_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_68_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_68_io_data_1_in_valid),
    .io_data_1_in_bits(PE_68_io_data_1_in_bits),
    .io_data_1_out_valid(PE_68_io_data_1_out_valid),
    .io_data_1_out_bits(PE_68_io_data_1_out_bits),
    .io_data_0_in_valid(PE_68_io_data_0_in_valid),
    .io_data_0_in_bits(PE_68_io_data_0_in_bits),
    .io_data_0_out_valid(PE_68_io_data_0_out_valid),
    .io_data_0_out_bits(PE_68_io_data_0_out_bits)
  );
  PE PE_69 ( // @[pe.scala 187:13]
    .clock(PE_69_clock),
    .reset(PE_69_reset),
    .io_data_2_out_valid(PE_69_io_data_2_out_valid),
    .io_data_2_out_bits(PE_69_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_69_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_69_io_data_1_in_valid),
    .io_data_1_in_bits(PE_69_io_data_1_in_bits),
    .io_data_1_out_valid(PE_69_io_data_1_out_valid),
    .io_data_1_out_bits(PE_69_io_data_1_out_bits),
    .io_data_0_in_valid(PE_69_io_data_0_in_valid),
    .io_data_0_in_bits(PE_69_io_data_0_in_bits),
    .io_data_0_out_valid(PE_69_io_data_0_out_valid),
    .io_data_0_out_bits(PE_69_io_data_0_out_bits)
  );
  PE PE_70 ( // @[pe.scala 187:13]
    .clock(PE_70_clock),
    .reset(PE_70_reset),
    .io_data_2_out_valid(PE_70_io_data_2_out_valid),
    .io_data_2_out_bits(PE_70_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_70_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_70_io_data_1_in_valid),
    .io_data_1_in_bits(PE_70_io_data_1_in_bits),
    .io_data_1_out_valid(PE_70_io_data_1_out_valid),
    .io_data_1_out_bits(PE_70_io_data_1_out_bits),
    .io_data_0_in_valid(PE_70_io_data_0_in_valid),
    .io_data_0_in_bits(PE_70_io_data_0_in_bits),
    .io_data_0_out_valid(PE_70_io_data_0_out_valid),
    .io_data_0_out_bits(PE_70_io_data_0_out_bits)
  );
  PE PE_71 ( // @[pe.scala 187:13]
    .clock(PE_71_clock),
    .reset(PE_71_reset),
    .io_data_2_out_valid(PE_71_io_data_2_out_valid),
    .io_data_2_out_bits(PE_71_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_71_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_71_io_data_1_in_valid),
    .io_data_1_in_bits(PE_71_io_data_1_in_bits),
    .io_data_1_out_valid(PE_71_io_data_1_out_valid),
    .io_data_1_out_bits(PE_71_io_data_1_out_bits),
    .io_data_0_in_valid(PE_71_io_data_0_in_valid),
    .io_data_0_in_bits(PE_71_io_data_0_in_bits),
    .io_data_0_out_valid(PE_71_io_data_0_out_valid),
    .io_data_0_out_bits(PE_71_io_data_0_out_bits)
  );
  PE PE_72 ( // @[pe.scala 187:13]
    .clock(PE_72_clock),
    .reset(PE_72_reset),
    .io_data_2_out_valid(PE_72_io_data_2_out_valid),
    .io_data_2_out_bits(PE_72_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_72_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_72_io_data_1_in_valid),
    .io_data_1_in_bits(PE_72_io_data_1_in_bits),
    .io_data_1_out_valid(PE_72_io_data_1_out_valid),
    .io_data_1_out_bits(PE_72_io_data_1_out_bits),
    .io_data_0_in_valid(PE_72_io_data_0_in_valid),
    .io_data_0_in_bits(PE_72_io_data_0_in_bits),
    .io_data_0_out_valid(PE_72_io_data_0_out_valid),
    .io_data_0_out_bits(PE_72_io_data_0_out_bits)
  );
  PE PE_73 ( // @[pe.scala 187:13]
    .clock(PE_73_clock),
    .reset(PE_73_reset),
    .io_data_2_out_valid(PE_73_io_data_2_out_valid),
    .io_data_2_out_bits(PE_73_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_73_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_73_io_data_1_in_valid),
    .io_data_1_in_bits(PE_73_io_data_1_in_bits),
    .io_data_1_out_valid(PE_73_io_data_1_out_valid),
    .io_data_1_out_bits(PE_73_io_data_1_out_bits),
    .io_data_0_in_valid(PE_73_io_data_0_in_valid),
    .io_data_0_in_bits(PE_73_io_data_0_in_bits),
    .io_data_0_out_valid(PE_73_io_data_0_out_valid),
    .io_data_0_out_bits(PE_73_io_data_0_out_bits)
  );
  PE PE_74 ( // @[pe.scala 187:13]
    .clock(PE_74_clock),
    .reset(PE_74_reset),
    .io_data_2_out_valid(PE_74_io_data_2_out_valid),
    .io_data_2_out_bits(PE_74_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_74_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_74_io_data_1_in_valid),
    .io_data_1_in_bits(PE_74_io_data_1_in_bits),
    .io_data_1_out_valid(PE_74_io_data_1_out_valid),
    .io_data_1_out_bits(PE_74_io_data_1_out_bits),
    .io_data_0_in_valid(PE_74_io_data_0_in_valid),
    .io_data_0_in_bits(PE_74_io_data_0_in_bits),
    .io_data_0_out_valid(PE_74_io_data_0_out_valid),
    .io_data_0_out_bits(PE_74_io_data_0_out_bits)
  );
  PE PE_75 ( // @[pe.scala 187:13]
    .clock(PE_75_clock),
    .reset(PE_75_reset),
    .io_data_2_out_valid(PE_75_io_data_2_out_valid),
    .io_data_2_out_bits(PE_75_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_75_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_75_io_data_1_in_valid),
    .io_data_1_in_bits(PE_75_io_data_1_in_bits),
    .io_data_1_out_valid(PE_75_io_data_1_out_valid),
    .io_data_1_out_bits(PE_75_io_data_1_out_bits),
    .io_data_0_in_valid(PE_75_io_data_0_in_valid),
    .io_data_0_in_bits(PE_75_io_data_0_in_bits),
    .io_data_0_out_valid(PE_75_io_data_0_out_valid),
    .io_data_0_out_bits(PE_75_io_data_0_out_bits)
  );
  PE PE_76 ( // @[pe.scala 187:13]
    .clock(PE_76_clock),
    .reset(PE_76_reset),
    .io_data_2_out_valid(PE_76_io_data_2_out_valid),
    .io_data_2_out_bits(PE_76_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_76_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_76_io_data_1_in_valid),
    .io_data_1_in_bits(PE_76_io_data_1_in_bits),
    .io_data_1_out_valid(PE_76_io_data_1_out_valid),
    .io_data_1_out_bits(PE_76_io_data_1_out_bits),
    .io_data_0_in_valid(PE_76_io_data_0_in_valid),
    .io_data_0_in_bits(PE_76_io_data_0_in_bits),
    .io_data_0_out_valid(PE_76_io_data_0_out_valid),
    .io_data_0_out_bits(PE_76_io_data_0_out_bits)
  );
  PE PE_77 ( // @[pe.scala 187:13]
    .clock(PE_77_clock),
    .reset(PE_77_reset),
    .io_data_2_out_valid(PE_77_io_data_2_out_valid),
    .io_data_2_out_bits(PE_77_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_77_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_77_io_data_1_in_valid),
    .io_data_1_in_bits(PE_77_io_data_1_in_bits),
    .io_data_1_out_valid(PE_77_io_data_1_out_valid),
    .io_data_1_out_bits(PE_77_io_data_1_out_bits),
    .io_data_0_in_valid(PE_77_io_data_0_in_valid),
    .io_data_0_in_bits(PE_77_io_data_0_in_bits),
    .io_data_0_out_valid(PE_77_io_data_0_out_valid),
    .io_data_0_out_bits(PE_77_io_data_0_out_bits)
  );
  PE PE_78 ( // @[pe.scala 187:13]
    .clock(PE_78_clock),
    .reset(PE_78_reset),
    .io_data_2_out_valid(PE_78_io_data_2_out_valid),
    .io_data_2_out_bits(PE_78_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_78_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_78_io_data_1_in_valid),
    .io_data_1_in_bits(PE_78_io_data_1_in_bits),
    .io_data_1_out_valid(PE_78_io_data_1_out_valid),
    .io_data_1_out_bits(PE_78_io_data_1_out_bits),
    .io_data_0_in_valid(PE_78_io_data_0_in_valid),
    .io_data_0_in_bits(PE_78_io_data_0_in_bits),
    .io_data_0_out_valid(PE_78_io_data_0_out_valid),
    .io_data_0_out_bits(PE_78_io_data_0_out_bits)
  );
  PE PE_79 ( // @[pe.scala 187:13]
    .clock(PE_79_clock),
    .reset(PE_79_reset),
    .io_data_2_out_valid(PE_79_io_data_2_out_valid),
    .io_data_2_out_bits(PE_79_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_79_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_79_io_data_1_in_valid),
    .io_data_1_in_bits(PE_79_io_data_1_in_bits),
    .io_data_1_out_valid(PE_79_io_data_1_out_valid),
    .io_data_1_out_bits(PE_79_io_data_1_out_bits),
    .io_data_0_in_valid(PE_79_io_data_0_in_valid),
    .io_data_0_in_bits(PE_79_io_data_0_in_bits),
    .io_data_0_out_valid(PE_79_io_data_0_out_valid),
    .io_data_0_out_bits(PE_79_io_data_0_out_bits)
  );
  PE PE_80 ( // @[pe.scala 187:13]
    .clock(PE_80_clock),
    .reset(PE_80_reset),
    .io_data_2_out_valid(PE_80_io_data_2_out_valid),
    .io_data_2_out_bits(PE_80_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_80_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_80_io_data_1_in_valid),
    .io_data_1_in_bits(PE_80_io_data_1_in_bits),
    .io_data_1_out_valid(PE_80_io_data_1_out_valid),
    .io_data_1_out_bits(PE_80_io_data_1_out_bits),
    .io_data_0_in_valid(PE_80_io_data_0_in_valid),
    .io_data_0_in_bits(PE_80_io_data_0_in_bits),
    .io_data_0_out_valid(PE_80_io_data_0_out_valid),
    .io_data_0_out_bits(PE_80_io_data_0_out_bits)
  );
  PE PE_81 ( // @[pe.scala 187:13]
    .clock(PE_81_clock),
    .reset(PE_81_reset),
    .io_data_2_out_valid(PE_81_io_data_2_out_valid),
    .io_data_2_out_bits(PE_81_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_81_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_81_io_data_1_in_valid),
    .io_data_1_in_bits(PE_81_io_data_1_in_bits),
    .io_data_1_out_valid(PE_81_io_data_1_out_valid),
    .io_data_1_out_bits(PE_81_io_data_1_out_bits),
    .io_data_0_in_valid(PE_81_io_data_0_in_valid),
    .io_data_0_in_bits(PE_81_io_data_0_in_bits),
    .io_data_0_out_valid(PE_81_io_data_0_out_valid),
    .io_data_0_out_bits(PE_81_io_data_0_out_bits)
  );
  PE PE_82 ( // @[pe.scala 187:13]
    .clock(PE_82_clock),
    .reset(PE_82_reset),
    .io_data_2_out_valid(PE_82_io_data_2_out_valid),
    .io_data_2_out_bits(PE_82_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_82_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_82_io_data_1_in_valid),
    .io_data_1_in_bits(PE_82_io_data_1_in_bits),
    .io_data_1_out_valid(PE_82_io_data_1_out_valid),
    .io_data_1_out_bits(PE_82_io_data_1_out_bits),
    .io_data_0_in_valid(PE_82_io_data_0_in_valid),
    .io_data_0_in_bits(PE_82_io_data_0_in_bits),
    .io_data_0_out_valid(PE_82_io_data_0_out_valid),
    .io_data_0_out_bits(PE_82_io_data_0_out_bits)
  );
  PE PE_83 ( // @[pe.scala 187:13]
    .clock(PE_83_clock),
    .reset(PE_83_reset),
    .io_data_2_out_valid(PE_83_io_data_2_out_valid),
    .io_data_2_out_bits(PE_83_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_83_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_83_io_data_1_in_valid),
    .io_data_1_in_bits(PE_83_io_data_1_in_bits),
    .io_data_1_out_valid(PE_83_io_data_1_out_valid),
    .io_data_1_out_bits(PE_83_io_data_1_out_bits),
    .io_data_0_in_valid(PE_83_io_data_0_in_valid),
    .io_data_0_in_bits(PE_83_io_data_0_in_bits),
    .io_data_0_out_valid(PE_83_io_data_0_out_valid),
    .io_data_0_out_bits(PE_83_io_data_0_out_bits)
  );
  PE PE_84 ( // @[pe.scala 187:13]
    .clock(PE_84_clock),
    .reset(PE_84_reset),
    .io_data_2_out_valid(PE_84_io_data_2_out_valid),
    .io_data_2_out_bits(PE_84_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_84_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_84_io_data_1_in_valid),
    .io_data_1_in_bits(PE_84_io_data_1_in_bits),
    .io_data_1_out_valid(PE_84_io_data_1_out_valid),
    .io_data_1_out_bits(PE_84_io_data_1_out_bits),
    .io_data_0_in_valid(PE_84_io_data_0_in_valid),
    .io_data_0_in_bits(PE_84_io_data_0_in_bits),
    .io_data_0_out_valid(PE_84_io_data_0_out_valid),
    .io_data_0_out_bits(PE_84_io_data_0_out_bits)
  );
  PE PE_85 ( // @[pe.scala 187:13]
    .clock(PE_85_clock),
    .reset(PE_85_reset),
    .io_data_2_out_valid(PE_85_io_data_2_out_valid),
    .io_data_2_out_bits(PE_85_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_85_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_85_io_data_1_in_valid),
    .io_data_1_in_bits(PE_85_io_data_1_in_bits),
    .io_data_1_out_valid(PE_85_io_data_1_out_valid),
    .io_data_1_out_bits(PE_85_io_data_1_out_bits),
    .io_data_0_in_valid(PE_85_io_data_0_in_valid),
    .io_data_0_in_bits(PE_85_io_data_0_in_bits),
    .io_data_0_out_valid(PE_85_io_data_0_out_valid),
    .io_data_0_out_bits(PE_85_io_data_0_out_bits)
  );
  PE PE_86 ( // @[pe.scala 187:13]
    .clock(PE_86_clock),
    .reset(PE_86_reset),
    .io_data_2_out_valid(PE_86_io_data_2_out_valid),
    .io_data_2_out_bits(PE_86_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_86_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_86_io_data_1_in_valid),
    .io_data_1_in_bits(PE_86_io_data_1_in_bits),
    .io_data_1_out_valid(PE_86_io_data_1_out_valid),
    .io_data_1_out_bits(PE_86_io_data_1_out_bits),
    .io_data_0_in_valid(PE_86_io_data_0_in_valid),
    .io_data_0_in_bits(PE_86_io_data_0_in_bits),
    .io_data_0_out_valid(PE_86_io_data_0_out_valid),
    .io_data_0_out_bits(PE_86_io_data_0_out_bits)
  );
  PE PE_87 ( // @[pe.scala 187:13]
    .clock(PE_87_clock),
    .reset(PE_87_reset),
    .io_data_2_out_valid(PE_87_io_data_2_out_valid),
    .io_data_2_out_bits(PE_87_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_87_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_87_io_data_1_in_valid),
    .io_data_1_in_bits(PE_87_io_data_1_in_bits),
    .io_data_1_out_valid(PE_87_io_data_1_out_valid),
    .io_data_1_out_bits(PE_87_io_data_1_out_bits),
    .io_data_0_in_valid(PE_87_io_data_0_in_valid),
    .io_data_0_in_bits(PE_87_io_data_0_in_bits),
    .io_data_0_out_valid(PE_87_io_data_0_out_valid),
    .io_data_0_out_bits(PE_87_io_data_0_out_bits)
  );
  PE PE_88 ( // @[pe.scala 187:13]
    .clock(PE_88_clock),
    .reset(PE_88_reset),
    .io_data_2_out_valid(PE_88_io_data_2_out_valid),
    .io_data_2_out_bits(PE_88_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_88_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_88_io_data_1_in_valid),
    .io_data_1_in_bits(PE_88_io_data_1_in_bits),
    .io_data_1_out_valid(PE_88_io_data_1_out_valid),
    .io_data_1_out_bits(PE_88_io_data_1_out_bits),
    .io_data_0_in_valid(PE_88_io_data_0_in_valid),
    .io_data_0_in_bits(PE_88_io_data_0_in_bits),
    .io_data_0_out_valid(PE_88_io_data_0_out_valid),
    .io_data_0_out_bits(PE_88_io_data_0_out_bits)
  );
  PE PE_89 ( // @[pe.scala 187:13]
    .clock(PE_89_clock),
    .reset(PE_89_reset),
    .io_data_2_out_valid(PE_89_io_data_2_out_valid),
    .io_data_2_out_bits(PE_89_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_89_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_89_io_data_1_in_valid),
    .io_data_1_in_bits(PE_89_io_data_1_in_bits),
    .io_data_1_out_valid(PE_89_io_data_1_out_valid),
    .io_data_1_out_bits(PE_89_io_data_1_out_bits),
    .io_data_0_in_valid(PE_89_io_data_0_in_valid),
    .io_data_0_in_bits(PE_89_io_data_0_in_bits),
    .io_data_0_out_valid(PE_89_io_data_0_out_valid),
    .io_data_0_out_bits(PE_89_io_data_0_out_bits)
  );
  PE PE_90 ( // @[pe.scala 187:13]
    .clock(PE_90_clock),
    .reset(PE_90_reset),
    .io_data_2_out_valid(PE_90_io_data_2_out_valid),
    .io_data_2_out_bits(PE_90_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_90_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_90_io_data_1_in_valid),
    .io_data_1_in_bits(PE_90_io_data_1_in_bits),
    .io_data_1_out_valid(PE_90_io_data_1_out_valid),
    .io_data_1_out_bits(PE_90_io_data_1_out_bits),
    .io_data_0_in_valid(PE_90_io_data_0_in_valid),
    .io_data_0_in_bits(PE_90_io_data_0_in_bits),
    .io_data_0_out_valid(PE_90_io_data_0_out_valid),
    .io_data_0_out_bits(PE_90_io_data_0_out_bits)
  );
  PE PE_91 ( // @[pe.scala 187:13]
    .clock(PE_91_clock),
    .reset(PE_91_reset),
    .io_data_2_out_valid(PE_91_io_data_2_out_valid),
    .io_data_2_out_bits(PE_91_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_91_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_91_io_data_1_in_valid),
    .io_data_1_in_bits(PE_91_io_data_1_in_bits),
    .io_data_1_out_valid(PE_91_io_data_1_out_valid),
    .io_data_1_out_bits(PE_91_io_data_1_out_bits),
    .io_data_0_in_valid(PE_91_io_data_0_in_valid),
    .io_data_0_in_bits(PE_91_io_data_0_in_bits),
    .io_data_0_out_valid(PE_91_io_data_0_out_valid),
    .io_data_0_out_bits(PE_91_io_data_0_out_bits)
  );
  PE PE_92 ( // @[pe.scala 187:13]
    .clock(PE_92_clock),
    .reset(PE_92_reset),
    .io_data_2_out_valid(PE_92_io_data_2_out_valid),
    .io_data_2_out_bits(PE_92_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_92_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_92_io_data_1_in_valid),
    .io_data_1_in_bits(PE_92_io_data_1_in_bits),
    .io_data_1_out_valid(PE_92_io_data_1_out_valid),
    .io_data_1_out_bits(PE_92_io_data_1_out_bits),
    .io_data_0_in_valid(PE_92_io_data_0_in_valid),
    .io_data_0_in_bits(PE_92_io_data_0_in_bits),
    .io_data_0_out_valid(PE_92_io_data_0_out_valid),
    .io_data_0_out_bits(PE_92_io_data_0_out_bits)
  );
  PE PE_93 ( // @[pe.scala 187:13]
    .clock(PE_93_clock),
    .reset(PE_93_reset),
    .io_data_2_out_valid(PE_93_io_data_2_out_valid),
    .io_data_2_out_bits(PE_93_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_93_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_93_io_data_1_in_valid),
    .io_data_1_in_bits(PE_93_io_data_1_in_bits),
    .io_data_1_out_valid(PE_93_io_data_1_out_valid),
    .io_data_1_out_bits(PE_93_io_data_1_out_bits),
    .io_data_0_in_valid(PE_93_io_data_0_in_valid),
    .io_data_0_in_bits(PE_93_io_data_0_in_bits),
    .io_data_0_out_valid(PE_93_io_data_0_out_valid),
    .io_data_0_out_bits(PE_93_io_data_0_out_bits)
  );
  PE PE_94 ( // @[pe.scala 187:13]
    .clock(PE_94_clock),
    .reset(PE_94_reset),
    .io_data_2_out_valid(PE_94_io_data_2_out_valid),
    .io_data_2_out_bits(PE_94_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_94_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_94_io_data_1_in_valid),
    .io_data_1_in_bits(PE_94_io_data_1_in_bits),
    .io_data_1_out_valid(PE_94_io_data_1_out_valid),
    .io_data_1_out_bits(PE_94_io_data_1_out_bits),
    .io_data_0_in_valid(PE_94_io_data_0_in_valid),
    .io_data_0_in_bits(PE_94_io_data_0_in_bits),
    .io_data_0_out_valid(PE_94_io_data_0_out_valid),
    .io_data_0_out_bits(PE_94_io_data_0_out_bits)
  );
  PE PE_95 ( // @[pe.scala 187:13]
    .clock(PE_95_clock),
    .reset(PE_95_reset),
    .io_data_2_out_valid(PE_95_io_data_2_out_valid),
    .io_data_2_out_bits(PE_95_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_95_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_95_io_data_1_in_valid),
    .io_data_1_in_bits(PE_95_io_data_1_in_bits),
    .io_data_1_out_valid(PE_95_io_data_1_out_valid),
    .io_data_1_out_bits(PE_95_io_data_1_out_bits),
    .io_data_0_in_valid(PE_95_io_data_0_in_valid),
    .io_data_0_in_bits(PE_95_io_data_0_in_bits),
    .io_data_0_out_valid(PE_95_io_data_0_out_valid),
    .io_data_0_out_bits(PE_95_io_data_0_out_bits)
  );
  PE PE_96 ( // @[pe.scala 187:13]
    .clock(PE_96_clock),
    .reset(PE_96_reset),
    .io_data_2_out_valid(PE_96_io_data_2_out_valid),
    .io_data_2_out_bits(PE_96_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_96_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_96_io_data_1_in_valid),
    .io_data_1_in_bits(PE_96_io_data_1_in_bits),
    .io_data_1_out_valid(PE_96_io_data_1_out_valid),
    .io_data_1_out_bits(PE_96_io_data_1_out_bits),
    .io_data_0_in_valid(PE_96_io_data_0_in_valid),
    .io_data_0_in_bits(PE_96_io_data_0_in_bits),
    .io_data_0_out_valid(PE_96_io_data_0_out_valid),
    .io_data_0_out_bits(PE_96_io_data_0_out_bits)
  );
  PE PE_97 ( // @[pe.scala 187:13]
    .clock(PE_97_clock),
    .reset(PE_97_reset),
    .io_data_2_out_valid(PE_97_io_data_2_out_valid),
    .io_data_2_out_bits(PE_97_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_97_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_97_io_data_1_in_valid),
    .io_data_1_in_bits(PE_97_io_data_1_in_bits),
    .io_data_1_out_valid(PE_97_io_data_1_out_valid),
    .io_data_1_out_bits(PE_97_io_data_1_out_bits),
    .io_data_0_in_valid(PE_97_io_data_0_in_valid),
    .io_data_0_in_bits(PE_97_io_data_0_in_bits),
    .io_data_0_out_valid(PE_97_io_data_0_out_valid),
    .io_data_0_out_bits(PE_97_io_data_0_out_bits)
  );
  PE PE_98 ( // @[pe.scala 187:13]
    .clock(PE_98_clock),
    .reset(PE_98_reset),
    .io_data_2_out_valid(PE_98_io_data_2_out_valid),
    .io_data_2_out_bits(PE_98_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_98_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_98_io_data_1_in_valid),
    .io_data_1_in_bits(PE_98_io_data_1_in_bits),
    .io_data_1_out_valid(PE_98_io_data_1_out_valid),
    .io_data_1_out_bits(PE_98_io_data_1_out_bits),
    .io_data_0_in_valid(PE_98_io_data_0_in_valid),
    .io_data_0_in_bits(PE_98_io_data_0_in_bits),
    .io_data_0_out_valid(PE_98_io_data_0_out_valid),
    .io_data_0_out_bits(PE_98_io_data_0_out_bits)
  );
  PE PE_99 ( // @[pe.scala 187:13]
    .clock(PE_99_clock),
    .reset(PE_99_reset),
    .io_data_2_out_valid(PE_99_io_data_2_out_valid),
    .io_data_2_out_bits(PE_99_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_99_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_99_io_data_1_in_valid),
    .io_data_1_in_bits(PE_99_io_data_1_in_bits),
    .io_data_1_out_valid(PE_99_io_data_1_out_valid),
    .io_data_1_out_bits(PE_99_io_data_1_out_bits),
    .io_data_0_in_valid(PE_99_io_data_0_in_valid),
    .io_data_0_in_bits(PE_99_io_data_0_in_bits),
    .io_data_0_out_valid(PE_99_io_data_0_out_valid),
    .io_data_0_out_bits(PE_99_io_data_0_out_bits)
  );
  PE PE_100 ( // @[pe.scala 187:13]
    .clock(PE_100_clock),
    .reset(PE_100_reset),
    .io_data_2_out_valid(PE_100_io_data_2_out_valid),
    .io_data_2_out_bits(PE_100_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_100_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_100_io_data_1_in_valid),
    .io_data_1_in_bits(PE_100_io_data_1_in_bits),
    .io_data_1_out_valid(PE_100_io_data_1_out_valid),
    .io_data_1_out_bits(PE_100_io_data_1_out_bits),
    .io_data_0_in_valid(PE_100_io_data_0_in_valid),
    .io_data_0_in_bits(PE_100_io_data_0_in_bits),
    .io_data_0_out_valid(PE_100_io_data_0_out_valid),
    .io_data_0_out_bits(PE_100_io_data_0_out_bits)
  );
  PE PE_101 ( // @[pe.scala 187:13]
    .clock(PE_101_clock),
    .reset(PE_101_reset),
    .io_data_2_out_valid(PE_101_io_data_2_out_valid),
    .io_data_2_out_bits(PE_101_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_101_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_101_io_data_1_in_valid),
    .io_data_1_in_bits(PE_101_io_data_1_in_bits),
    .io_data_1_out_valid(PE_101_io_data_1_out_valid),
    .io_data_1_out_bits(PE_101_io_data_1_out_bits),
    .io_data_0_in_valid(PE_101_io_data_0_in_valid),
    .io_data_0_in_bits(PE_101_io_data_0_in_bits),
    .io_data_0_out_valid(PE_101_io_data_0_out_valid),
    .io_data_0_out_bits(PE_101_io_data_0_out_bits)
  );
  PE PE_102 ( // @[pe.scala 187:13]
    .clock(PE_102_clock),
    .reset(PE_102_reset),
    .io_data_2_out_valid(PE_102_io_data_2_out_valid),
    .io_data_2_out_bits(PE_102_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_102_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_102_io_data_1_in_valid),
    .io_data_1_in_bits(PE_102_io_data_1_in_bits),
    .io_data_1_out_valid(PE_102_io_data_1_out_valid),
    .io_data_1_out_bits(PE_102_io_data_1_out_bits),
    .io_data_0_in_valid(PE_102_io_data_0_in_valid),
    .io_data_0_in_bits(PE_102_io_data_0_in_bits),
    .io_data_0_out_valid(PE_102_io_data_0_out_valid),
    .io_data_0_out_bits(PE_102_io_data_0_out_bits)
  );
  PE PE_103 ( // @[pe.scala 187:13]
    .clock(PE_103_clock),
    .reset(PE_103_reset),
    .io_data_2_out_valid(PE_103_io_data_2_out_valid),
    .io_data_2_out_bits(PE_103_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_103_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_103_io_data_1_in_valid),
    .io_data_1_in_bits(PE_103_io_data_1_in_bits),
    .io_data_1_out_valid(PE_103_io_data_1_out_valid),
    .io_data_1_out_bits(PE_103_io_data_1_out_bits),
    .io_data_0_in_valid(PE_103_io_data_0_in_valid),
    .io_data_0_in_bits(PE_103_io_data_0_in_bits),
    .io_data_0_out_valid(PE_103_io_data_0_out_valid),
    .io_data_0_out_bits(PE_103_io_data_0_out_bits)
  );
  PE PE_104 ( // @[pe.scala 187:13]
    .clock(PE_104_clock),
    .reset(PE_104_reset),
    .io_data_2_out_valid(PE_104_io_data_2_out_valid),
    .io_data_2_out_bits(PE_104_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_104_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_104_io_data_1_in_valid),
    .io_data_1_in_bits(PE_104_io_data_1_in_bits),
    .io_data_1_out_valid(PE_104_io_data_1_out_valid),
    .io_data_1_out_bits(PE_104_io_data_1_out_bits),
    .io_data_0_in_valid(PE_104_io_data_0_in_valid),
    .io_data_0_in_bits(PE_104_io_data_0_in_bits),
    .io_data_0_out_valid(PE_104_io_data_0_out_valid),
    .io_data_0_out_bits(PE_104_io_data_0_out_bits)
  );
  PE PE_105 ( // @[pe.scala 187:13]
    .clock(PE_105_clock),
    .reset(PE_105_reset),
    .io_data_2_out_valid(PE_105_io_data_2_out_valid),
    .io_data_2_out_bits(PE_105_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_105_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_105_io_data_1_in_valid),
    .io_data_1_in_bits(PE_105_io_data_1_in_bits),
    .io_data_1_out_valid(PE_105_io_data_1_out_valid),
    .io_data_1_out_bits(PE_105_io_data_1_out_bits),
    .io_data_0_in_valid(PE_105_io_data_0_in_valid),
    .io_data_0_in_bits(PE_105_io_data_0_in_bits),
    .io_data_0_out_valid(PE_105_io_data_0_out_valid),
    .io_data_0_out_bits(PE_105_io_data_0_out_bits)
  );
  PE PE_106 ( // @[pe.scala 187:13]
    .clock(PE_106_clock),
    .reset(PE_106_reset),
    .io_data_2_out_valid(PE_106_io_data_2_out_valid),
    .io_data_2_out_bits(PE_106_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_106_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_106_io_data_1_in_valid),
    .io_data_1_in_bits(PE_106_io_data_1_in_bits),
    .io_data_1_out_valid(PE_106_io_data_1_out_valid),
    .io_data_1_out_bits(PE_106_io_data_1_out_bits),
    .io_data_0_in_valid(PE_106_io_data_0_in_valid),
    .io_data_0_in_bits(PE_106_io_data_0_in_bits),
    .io_data_0_out_valid(PE_106_io_data_0_out_valid),
    .io_data_0_out_bits(PE_106_io_data_0_out_bits)
  );
  PE PE_107 ( // @[pe.scala 187:13]
    .clock(PE_107_clock),
    .reset(PE_107_reset),
    .io_data_2_out_valid(PE_107_io_data_2_out_valid),
    .io_data_2_out_bits(PE_107_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_107_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_107_io_data_1_in_valid),
    .io_data_1_in_bits(PE_107_io_data_1_in_bits),
    .io_data_1_out_valid(PE_107_io_data_1_out_valid),
    .io_data_1_out_bits(PE_107_io_data_1_out_bits),
    .io_data_0_in_valid(PE_107_io_data_0_in_valid),
    .io_data_0_in_bits(PE_107_io_data_0_in_bits),
    .io_data_0_out_valid(PE_107_io_data_0_out_valid),
    .io_data_0_out_bits(PE_107_io_data_0_out_bits)
  );
  PE PE_108 ( // @[pe.scala 187:13]
    .clock(PE_108_clock),
    .reset(PE_108_reset),
    .io_data_2_out_valid(PE_108_io_data_2_out_valid),
    .io_data_2_out_bits(PE_108_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_108_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_108_io_data_1_in_valid),
    .io_data_1_in_bits(PE_108_io_data_1_in_bits),
    .io_data_1_out_valid(PE_108_io_data_1_out_valid),
    .io_data_1_out_bits(PE_108_io_data_1_out_bits),
    .io_data_0_in_valid(PE_108_io_data_0_in_valid),
    .io_data_0_in_bits(PE_108_io_data_0_in_bits),
    .io_data_0_out_valid(PE_108_io_data_0_out_valid),
    .io_data_0_out_bits(PE_108_io_data_0_out_bits)
  );
  PE PE_109 ( // @[pe.scala 187:13]
    .clock(PE_109_clock),
    .reset(PE_109_reset),
    .io_data_2_out_valid(PE_109_io_data_2_out_valid),
    .io_data_2_out_bits(PE_109_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_109_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_109_io_data_1_in_valid),
    .io_data_1_in_bits(PE_109_io_data_1_in_bits),
    .io_data_1_out_valid(PE_109_io_data_1_out_valid),
    .io_data_1_out_bits(PE_109_io_data_1_out_bits),
    .io_data_0_in_valid(PE_109_io_data_0_in_valid),
    .io_data_0_in_bits(PE_109_io_data_0_in_bits),
    .io_data_0_out_valid(PE_109_io_data_0_out_valid),
    .io_data_0_out_bits(PE_109_io_data_0_out_bits)
  );
  PE PE_110 ( // @[pe.scala 187:13]
    .clock(PE_110_clock),
    .reset(PE_110_reset),
    .io_data_2_out_valid(PE_110_io_data_2_out_valid),
    .io_data_2_out_bits(PE_110_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_110_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_110_io_data_1_in_valid),
    .io_data_1_in_bits(PE_110_io_data_1_in_bits),
    .io_data_1_out_valid(PE_110_io_data_1_out_valid),
    .io_data_1_out_bits(PE_110_io_data_1_out_bits),
    .io_data_0_in_valid(PE_110_io_data_0_in_valid),
    .io_data_0_in_bits(PE_110_io_data_0_in_bits),
    .io_data_0_out_valid(PE_110_io_data_0_out_valid),
    .io_data_0_out_bits(PE_110_io_data_0_out_bits)
  );
  PE PE_111 ( // @[pe.scala 187:13]
    .clock(PE_111_clock),
    .reset(PE_111_reset),
    .io_data_2_out_valid(PE_111_io_data_2_out_valid),
    .io_data_2_out_bits(PE_111_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_111_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_111_io_data_1_in_valid),
    .io_data_1_in_bits(PE_111_io_data_1_in_bits),
    .io_data_1_out_valid(PE_111_io_data_1_out_valid),
    .io_data_1_out_bits(PE_111_io_data_1_out_bits),
    .io_data_0_in_valid(PE_111_io_data_0_in_valid),
    .io_data_0_in_bits(PE_111_io_data_0_in_bits),
    .io_data_0_out_valid(PE_111_io_data_0_out_valid),
    .io_data_0_out_bits(PE_111_io_data_0_out_bits)
  );
  PE PE_112 ( // @[pe.scala 187:13]
    .clock(PE_112_clock),
    .reset(PE_112_reset),
    .io_data_2_out_valid(PE_112_io_data_2_out_valid),
    .io_data_2_out_bits(PE_112_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_112_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_112_io_data_1_in_valid),
    .io_data_1_in_bits(PE_112_io_data_1_in_bits),
    .io_data_1_out_valid(PE_112_io_data_1_out_valid),
    .io_data_1_out_bits(PE_112_io_data_1_out_bits),
    .io_data_0_in_valid(PE_112_io_data_0_in_valid),
    .io_data_0_in_bits(PE_112_io_data_0_in_bits),
    .io_data_0_out_valid(PE_112_io_data_0_out_valid),
    .io_data_0_out_bits(PE_112_io_data_0_out_bits)
  );
  PE PE_113 ( // @[pe.scala 187:13]
    .clock(PE_113_clock),
    .reset(PE_113_reset),
    .io_data_2_out_valid(PE_113_io_data_2_out_valid),
    .io_data_2_out_bits(PE_113_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_113_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_113_io_data_1_in_valid),
    .io_data_1_in_bits(PE_113_io_data_1_in_bits),
    .io_data_1_out_valid(PE_113_io_data_1_out_valid),
    .io_data_1_out_bits(PE_113_io_data_1_out_bits),
    .io_data_0_in_valid(PE_113_io_data_0_in_valid),
    .io_data_0_in_bits(PE_113_io_data_0_in_bits),
    .io_data_0_out_valid(PE_113_io_data_0_out_valid),
    .io_data_0_out_bits(PE_113_io_data_0_out_bits)
  );
  PE PE_114 ( // @[pe.scala 187:13]
    .clock(PE_114_clock),
    .reset(PE_114_reset),
    .io_data_2_out_valid(PE_114_io_data_2_out_valid),
    .io_data_2_out_bits(PE_114_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_114_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_114_io_data_1_in_valid),
    .io_data_1_in_bits(PE_114_io_data_1_in_bits),
    .io_data_1_out_valid(PE_114_io_data_1_out_valid),
    .io_data_1_out_bits(PE_114_io_data_1_out_bits),
    .io_data_0_in_valid(PE_114_io_data_0_in_valid),
    .io_data_0_in_bits(PE_114_io_data_0_in_bits),
    .io_data_0_out_valid(PE_114_io_data_0_out_valid),
    .io_data_0_out_bits(PE_114_io_data_0_out_bits)
  );
  PE PE_115 ( // @[pe.scala 187:13]
    .clock(PE_115_clock),
    .reset(PE_115_reset),
    .io_data_2_out_valid(PE_115_io_data_2_out_valid),
    .io_data_2_out_bits(PE_115_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_115_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_115_io_data_1_in_valid),
    .io_data_1_in_bits(PE_115_io_data_1_in_bits),
    .io_data_1_out_valid(PE_115_io_data_1_out_valid),
    .io_data_1_out_bits(PE_115_io_data_1_out_bits),
    .io_data_0_in_valid(PE_115_io_data_0_in_valid),
    .io_data_0_in_bits(PE_115_io_data_0_in_bits),
    .io_data_0_out_valid(PE_115_io_data_0_out_valid),
    .io_data_0_out_bits(PE_115_io_data_0_out_bits)
  );
  PE PE_116 ( // @[pe.scala 187:13]
    .clock(PE_116_clock),
    .reset(PE_116_reset),
    .io_data_2_out_valid(PE_116_io_data_2_out_valid),
    .io_data_2_out_bits(PE_116_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_116_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_116_io_data_1_in_valid),
    .io_data_1_in_bits(PE_116_io_data_1_in_bits),
    .io_data_1_out_valid(PE_116_io_data_1_out_valid),
    .io_data_1_out_bits(PE_116_io_data_1_out_bits),
    .io_data_0_in_valid(PE_116_io_data_0_in_valid),
    .io_data_0_in_bits(PE_116_io_data_0_in_bits),
    .io_data_0_out_valid(PE_116_io_data_0_out_valid),
    .io_data_0_out_bits(PE_116_io_data_0_out_bits)
  );
  PE PE_117 ( // @[pe.scala 187:13]
    .clock(PE_117_clock),
    .reset(PE_117_reset),
    .io_data_2_out_valid(PE_117_io_data_2_out_valid),
    .io_data_2_out_bits(PE_117_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_117_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_117_io_data_1_in_valid),
    .io_data_1_in_bits(PE_117_io_data_1_in_bits),
    .io_data_1_out_valid(PE_117_io_data_1_out_valid),
    .io_data_1_out_bits(PE_117_io_data_1_out_bits),
    .io_data_0_in_valid(PE_117_io_data_0_in_valid),
    .io_data_0_in_bits(PE_117_io_data_0_in_bits),
    .io_data_0_out_valid(PE_117_io_data_0_out_valid),
    .io_data_0_out_bits(PE_117_io_data_0_out_bits)
  );
  PE PE_118 ( // @[pe.scala 187:13]
    .clock(PE_118_clock),
    .reset(PE_118_reset),
    .io_data_2_out_valid(PE_118_io_data_2_out_valid),
    .io_data_2_out_bits(PE_118_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_118_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_118_io_data_1_in_valid),
    .io_data_1_in_bits(PE_118_io_data_1_in_bits),
    .io_data_1_out_valid(PE_118_io_data_1_out_valid),
    .io_data_1_out_bits(PE_118_io_data_1_out_bits),
    .io_data_0_in_valid(PE_118_io_data_0_in_valid),
    .io_data_0_in_bits(PE_118_io_data_0_in_bits),
    .io_data_0_out_valid(PE_118_io_data_0_out_valid),
    .io_data_0_out_bits(PE_118_io_data_0_out_bits)
  );
  PE PE_119 ( // @[pe.scala 187:13]
    .clock(PE_119_clock),
    .reset(PE_119_reset),
    .io_data_2_out_valid(PE_119_io_data_2_out_valid),
    .io_data_2_out_bits(PE_119_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_119_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_119_io_data_1_in_valid),
    .io_data_1_in_bits(PE_119_io_data_1_in_bits),
    .io_data_1_out_valid(PE_119_io_data_1_out_valid),
    .io_data_1_out_bits(PE_119_io_data_1_out_bits),
    .io_data_0_in_valid(PE_119_io_data_0_in_valid),
    .io_data_0_in_bits(PE_119_io_data_0_in_bits),
    .io_data_0_out_valid(PE_119_io_data_0_out_valid),
    .io_data_0_out_bits(PE_119_io_data_0_out_bits)
  );
  PE PE_120 ( // @[pe.scala 187:13]
    .clock(PE_120_clock),
    .reset(PE_120_reset),
    .io_data_2_out_valid(PE_120_io_data_2_out_valid),
    .io_data_2_out_bits(PE_120_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_120_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_120_io_data_1_in_valid),
    .io_data_1_in_bits(PE_120_io_data_1_in_bits),
    .io_data_1_out_valid(PE_120_io_data_1_out_valid),
    .io_data_1_out_bits(PE_120_io_data_1_out_bits),
    .io_data_0_in_valid(PE_120_io_data_0_in_valid),
    .io_data_0_in_bits(PE_120_io_data_0_in_bits),
    .io_data_0_out_valid(PE_120_io_data_0_out_valid),
    .io_data_0_out_bits(PE_120_io_data_0_out_bits)
  );
  PE PE_121 ( // @[pe.scala 187:13]
    .clock(PE_121_clock),
    .reset(PE_121_reset),
    .io_data_2_out_valid(PE_121_io_data_2_out_valid),
    .io_data_2_out_bits(PE_121_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_121_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_121_io_data_1_in_valid),
    .io_data_1_in_bits(PE_121_io_data_1_in_bits),
    .io_data_1_out_valid(PE_121_io_data_1_out_valid),
    .io_data_1_out_bits(PE_121_io_data_1_out_bits),
    .io_data_0_in_valid(PE_121_io_data_0_in_valid),
    .io_data_0_in_bits(PE_121_io_data_0_in_bits),
    .io_data_0_out_valid(PE_121_io_data_0_out_valid),
    .io_data_0_out_bits(PE_121_io_data_0_out_bits)
  );
  PE PE_122 ( // @[pe.scala 187:13]
    .clock(PE_122_clock),
    .reset(PE_122_reset),
    .io_data_2_out_valid(PE_122_io_data_2_out_valid),
    .io_data_2_out_bits(PE_122_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_122_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_122_io_data_1_in_valid),
    .io_data_1_in_bits(PE_122_io_data_1_in_bits),
    .io_data_1_out_valid(PE_122_io_data_1_out_valid),
    .io_data_1_out_bits(PE_122_io_data_1_out_bits),
    .io_data_0_in_valid(PE_122_io_data_0_in_valid),
    .io_data_0_in_bits(PE_122_io_data_0_in_bits),
    .io_data_0_out_valid(PE_122_io_data_0_out_valid),
    .io_data_0_out_bits(PE_122_io_data_0_out_bits)
  );
  PE PE_123 ( // @[pe.scala 187:13]
    .clock(PE_123_clock),
    .reset(PE_123_reset),
    .io_data_2_out_valid(PE_123_io_data_2_out_valid),
    .io_data_2_out_bits(PE_123_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_123_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_123_io_data_1_in_valid),
    .io_data_1_in_bits(PE_123_io_data_1_in_bits),
    .io_data_1_out_valid(PE_123_io_data_1_out_valid),
    .io_data_1_out_bits(PE_123_io_data_1_out_bits),
    .io_data_0_in_valid(PE_123_io_data_0_in_valid),
    .io_data_0_in_bits(PE_123_io_data_0_in_bits),
    .io_data_0_out_valid(PE_123_io_data_0_out_valid),
    .io_data_0_out_bits(PE_123_io_data_0_out_bits)
  );
  PE PE_124 ( // @[pe.scala 187:13]
    .clock(PE_124_clock),
    .reset(PE_124_reset),
    .io_data_2_out_valid(PE_124_io_data_2_out_valid),
    .io_data_2_out_bits(PE_124_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_124_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_124_io_data_1_in_valid),
    .io_data_1_in_bits(PE_124_io_data_1_in_bits),
    .io_data_1_out_valid(PE_124_io_data_1_out_valid),
    .io_data_1_out_bits(PE_124_io_data_1_out_bits),
    .io_data_0_in_valid(PE_124_io_data_0_in_valid),
    .io_data_0_in_bits(PE_124_io_data_0_in_bits),
    .io_data_0_out_valid(PE_124_io_data_0_out_valid),
    .io_data_0_out_bits(PE_124_io_data_0_out_bits)
  );
  PE PE_125 ( // @[pe.scala 187:13]
    .clock(PE_125_clock),
    .reset(PE_125_reset),
    .io_data_2_out_valid(PE_125_io_data_2_out_valid),
    .io_data_2_out_bits(PE_125_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_125_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_125_io_data_1_in_valid),
    .io_data_1_in_bits(PE_125_io_data_1_in_bits),
    .io_data_1_out_valid(PE_125_io_data_1_out_valid),
    .io_data_1_out_bits(PE_125_io_data_1_out_bits),
    .io_data_0_in_valid(PE_125_io_data_0_in_valid),
    .io_data_0_in_bits(PE_125_io_data_0_in_bits),
    .io_data_0_out_valid(PE_125_io_data_0_out_valid),
    .io_data_0_out_bits(PE_125_io_data_0_out_bits)
  );
  PE PE_126 ( // @[pe.scala 187:13]
    .clock(PE_126_clock),
    .reset(PE_126_reset),
    .io_data_2_out_valid(PE_126_io_data_2_out_valid),
    .io_data_2_out_bits(PE_126_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_126_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_126_io_data_1_in_valid),
    .io_data_1_in_bits(PE_126_io_data_1_in_bits),
    .io_data_1_out_valid(PE_126_io_data_1_out_valid),
    .io_data_1_out_bits(PE_126_io_data_1_out_bits),
    .io_data_0_in_valid(PE_126_io_data_0_in_valid),
    .io_data_0_in_bits(PE_126_io_data_0_in_bits),
    .io_data_0_out_valid(PE_126_io_data_0_out_valid),
    .io_data_0_out_bits(PE_126_io_data_0_out_bits)
  );
  PE PE_127 ( // @[pe.scala 187:13]
    .clock(PE_127_clock),
    .reset(PE_127_reset),
    .io_data_2_out_valid(PE_127_io_data_2_out_valid),
    .io_data_2_out_bits(PE_127_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_127_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_127_io_data_1_in_valid),
    .io_data_1_in_bits(PE_127_io_data_1_in_bits),
    .io_data_1_out_valid(PE_127_io_data_1_out_valid),
    .io_data_1_out_bits(PE_127_io_data_1_out_bits),
    .io_data_0_in_valid(PE_127_io_data_0_in_valid),
    .io_data_0_in_bits(PE_127_io_data_0_in_bits),
    .io_data_0_out_valid(PE_127_io_data_0_out_valid),
    .io_data_0_out_bits(PE_127_io_data_0_out_bits)
  );
  PE PE_128 ( // @[pe.scala 187:13]
    .clock(PE_128_clock),
    .reset(PE_128_reset),
    .io_data_2_out_valid(PE_128_io_data_2_out_valid),
    .io_data_2_out_bits(PE_128_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_128_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_128_io_data_1_in_valid),
    .io_data_1_in_bits(PE_128_io_data_1_in_bits),
    .io_data_1_out_valid(PE_128_io_data_1_out_valid),
    .io_data_1_out_bits(PE_128_io_data_1_out_bits),
    .io_data_0_in_valid(PE_128_io_data_0_in_valid),
    .io_data_0_in_bits(PE_128_io_data_0_in_bits),
    .io_data_0_out_valid(PE_128_io_data_0_out_valid),
    .io_data_0_out_bits(PE_128_io_data_0_out_bits)
  );
  PE PE_129 ( // @[pe.scala 187:13]
    .clock(PE_129_clock),
    .reset(PE_129_reset),
    .io_data_2_out_valid(PE_129_io_data_2_out_valid),
    .io_data_2_out_bits(PE_129_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_129_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_129_io_data_1_in_valid),
    .io_data_1_in_bits(PE_129_io_data_1_in_bits),
    .io_data_1_out_valid(PE_129_io_data_1_out_valid),
    .io_data_1_out_bits(PE_129_io_data_1_out_bits),
    .io_data_0_in_valid(PE_129_io_data_0_in_valid),
    .io_data_0_in_bits(PE_129_io_data_0_in_bits),
    .io_data_0_out_valid(PE_129_io_data_0_out_valid),
    .io_data_0_out_bits(PE_129_io_data_0_out_bits)
  );
  PE PE_130 ( // @[pe.scala 187:13]
    .clock(PE_130_clock),
    .reset(PE_130_reset),
    .io_data_2_out_valid(PE_130_io_data_2_out_valid),
    .io_data_2_out_bits(PE_130_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_130_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_130_io_data_1_in_valid),
    .io_data_1_in_bits(PE_130_io_data_1_in_bits),
    .io_data_1_out_valid(PE_130_io_data_1_out_valid),
    .io_data_1_out_bits(PE_130_io_data_1_out_bits),
    .io_data_0_in_valid(PE_130_io_data_0_in_valid),
    .io_data_0_in_bits(PE_130_io_data_0_in_bits),
    .io_data_0_out_valid(PE_130_io_data_0_out_valid),
    .io_data_0_out_bits(PE_130_io_data_0_out_bits)
  );
  PE PE_131 ( // @[pe.scala 187:13]
    .clock(PE_131_clock),
    .reset(PE_131_reset),
    .io_data_2_out_valid(PE_131_io_data_2_out_valid),
    .io_data_2_out_bits(PE_131_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_131_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_131_io_data_1_in_valid),
    .io_data_1_in_bits(PE_131_io_data_1_in_bits),
    .io_data_1_out_valid(PE_131_io_data_1_out_valid),
    .io_data_1_out_bits(PE_131_io_data_1_out_bits),
    .io_data_0_in_valid(PE_131_io_data_0_in_valid),
    .io_data_0_in_bits(PE_131_io_data_0_in_bits),
    .io_data_0_out_valid(PE_131_io_data_0_out_valid),
    .io_data_0_out_bits(PE_131_io_data_0_out_bits)
  );
  PE PE_132 ( // @[pe.scala 187:13]
    .clock(PE_132_clock),
    .reset(PE_132_reset),
    .io_data_2_out_valid(PE_132_io_data_2_out_valid),
    .io_data_2_out_bits(PE_132_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_132_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_132_io_data_1_in_valid),
    .io_data_1_in_bits(PE_132_io_data_1_in_bits),
    .io_data_1_out_valid(PE_132_io_data_1_out_valid),
    .io_data_1_out_bits(PE_132_io_data_1_out_bits),
    .io_data_0_in_valid(PE_132_io_data_0_in_valid),
    .io_data_0_in_bits(PE_132_io_data_0_in_bits),
    .io_data_0_out_valid(PE_132_io_data_0_out_valid),
    .io_data_0_out_bits(PE_132_io_data_0_out_bits)
  );
  PE PE_133 ( // @[pe.scala 187:13]
    .clock(PE_133_clock),
    .reset(PE_133_reset),
    .io_data_2_out_valid(PE_133_io_data_2_out_valid),
    .io_data_2_out_bits(PE_133_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_133_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_133_io_data_1_in_valid),
    .io_data_1_in_bits(PE_133_io_data_1_in_bits),
    .io_data_1_out_valid(PE_133_io_data_1_out_valid),
    .io_data_1_out_bits(PE_133_io_data_1_out_bits),
    .io_data_0_in_valid(PE_133_io_data_0_in_valid),
    .io_data_0_in_bits(PE_133_io_data_0_in_bits),
    .io_data_0_out_valid(PE_133_io_data_0_out_valid),
    .io_data_0_out_bits(PE_133_io_data_0_out_bits)
  );
  PE PE_134 ( // @[pe.scala 187:13]
    .clock(PE_134_clock),
    .reset(PE_134_reset),
    .io_data_2_out_valid(PE_134_io_data_2_out_valid),
    .io_data_2_out_bits(PE_134_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_134_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_134_io_data_1_in_valid),
    .io_data_1_in_bits(PE_134_io_data_1_in_bits),
    .io_data_1_out_valid(PE_134_io_data_1_out_valid),
    .io_data_1_out_bits(PE_134_io_data_1_out_bits),
    .io_data_0_in_valid(PE_134_io_data_0_in_valid),
    .io_data_0_in_bits(PE_134_io_data_0_in_bits),
    .io_data_0_out_valid(PE_134_io_data_0_out_valid),
    .io_data_0_out_bits(PE_134_io_data_0_out_bits)
  );
  PE PE_135 ( // @[pe.scala 187:13]
    .clock(PE_135_clock),
    .reset(PE_135_reset),
    .io_data_2_out_valid(PE_135_io_data_2_out_valid),
    .io_data_2_out_bits(PE_135_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_135_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_135_io_data_1_in_valid),
    .io_data_1_in_bits(PE_135_io_data_1_in_bits),
    .io_data_1_out_valid(PE_135_io_data_1_out_valid),
    .io_data_1_out_bits(PE_135_io_data_1_out_bits),
    .io_data_0_in_valid(PE_135_io_data_0_in_valid),
    .io_data_0_in_bits(PE_135_io_data_0_in_bits),
    .io_data_0_out_valid(PE_135_io_data_0_out_valid),
    .io_data_0_out_bits(PE_135_io_data_0_out_bits)
  );
  PE PE_136 ( // @[pe.scala 187:13]
    .clock(PE_136_clock),
    .reset(PE_136_reset),
    .io_data_2_out_valid(PE_136_io_data_2_out_valid),
    .io_data_2_out_bits(PE_136_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_136_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_136_io_data_1_in_valid),
    .io_data_1_in_bits(PE_136_io_data_1_in_bits),
    .io_data_1_out_valid(PE_136_io_data_1_out_valid),
    .io_data_1_out_bits(PE_136_io_data_1_out_bits),
    .io_data_0_in_valid(PE_136_io_data_0_in_valid),
    .io_data_0_in_bits(PE_136_io_data_0_in_bits),
    .io_data_0_out_valid(PE_136_io_data_0_out_valid),
    .io_data_0_out_bits(PE_136_io_data_0_out_bits)
  );
  PE PE_137 ( // @[pe.scala 187:13]
    .clock(PE_137_clock),
    .reset(PE_137_reset),
    .io_data_2_out_valid(PE_137_io_data_2_out_valid),
    .io_data_2_out_bits(PE_137_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_137_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_137_io_data_1_in_valid),
    .io_data_1_in_bits(PE_137_io_data_1_in_bits),
    .io_data_1_out_valid(PE_137_io_data_1_out_valid),
    .io_data_1_out_bits(PE_137_io_data_1_out_bits),
    .io_data_0_in_valid(PE_137_io_data_0_in_valid),
    .io_data_0_in_bits(PE_137_io_data_0_in_bits),
    .io_data_0_out_valid(PE_137_io_data_0_out_valid),
    .io_data_0_out_bits(PE_137_io_data_0_out_bits)
  );
  PE PE_138 ( // @[pe.scala 187:13]
    .clock(PE_138_clock),
    .reset(PE_138_reset),
    .io_data_2_out_valid(PE_138_io_data_2_out_valid),
    .io_data_2_out_bits(PE_138_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_138_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_138_io_data_1_in_valid),
    .io_data_1_in_bits(PE_138_io_data_1_in_bits),
    .io_data_1_out_valid(PE_138_io_data_1_out_valid),
    .io_data_1_out_bits(PE_138_io_data_1_out_bits),
    .io_data_0_in_valid(PE_138_io_data_0_in_valid),
    .io_data_0_in_bits(PE_138_io_data_0_in_bits),
    .io_data_0_out_valid(PE_138_io_data_0_out_valid),
    .io_data_0_out_bits(PE_138_io_data_0_out_bits)
  );
  PE PE_139 ( // @[pe.scala 187:13]
    .clock(PE_139_clock),
    .reset(PE_139_reset),
    .io_data_2_out_valid(PE_139_io_data_2_out_valid),
    .io_data_2_out_bits(PE_139_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_139_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_139_io_data_1_in_valid),
    .io_data_1_in_bits(PE_139_io_data_1_in_bits),
    .io_data_1_out_valid(PE_139_io_data_1_out_valid),
    .io_data_1_out_bits(PE_139_io_data_1_out_bits),
    .io_data_0_in_valid(PE_139_io_data_0_in_valid),
    .io_data_0_in_bits(PE_139_io_data_0_in_bits),
    .io_data_0_out_valid(PE_139_io_data_0_out_valid),
    .io_data_0_out_bits(PE_139_io_data_0_out_bits)
  );
  PE PE_140 ( // @[pe.scala 187:13]
    .clock(PE_140_clock),
    .reset(PE_140_reset),
    .io_data_2_out_valid(PE_140_io_data_2_out_valid),
    .io_data_2_out_bits(PE_140_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_140_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_140_io_data_1_in_valid),
    .io_data_1_in_bits(PE_140_io_data_1_in_bits),
    .io_data_1_out_valid(PE_140_io_data_1_out_valid),
    .io_data_1_out_bits(PE_140_io_data_1_out_bits),
    .io_data_0_in_valid(PE_140_io_data_0_in_valid),
    .io_data_0_in_bits(PE_140_io_data_0_in_bits),
    .io_data_0_out_valid(PE_140_io_data_0_out_valid),
    .io_data_0_out_bits(PE_140_io_data_0_out_bits)
  );
  PE PE_141 ( // @[pe.scala 187:13]
    .clock(PE_141_clock),
    .reset(PE_141_reset),
    .io_data_2_out_valid(PE_141_io_data_2_out_valid),
    .io_data_2_out_bits(PE_141_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_141_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_141_io_data_1_in_valid),
    .io_data_1_in_bits(PE_141_io_data_1_in_bits),
    .io_data_1_out_valid(PE_141_io_data_1_out_valid),
    .io_data_1_out_bits(PE_141_io_data_1_out_bits),
    .io_data_0_in_valid(PE_141_io_data_0_in_valid),
    .io_data_0_in_bits(PE_141_io_data_0_in_bits),
    .io_data_0_out_valid(PE_141_io_data_0_out_valid),
    .io_data_0_out_bits(PE_141_io_data_0_out_bits)
  );
  PE PE_142 ( // @[pe.scala 187:13]
    .clock(PE_142_clock),
    .reset(PE_142_reset),
    .io_data_2_out_valid(PE_142_io_data_2_out_valid),
    .io_data_2_out_bits(PE_142_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_142_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_142_io_data_1_in_valid),
    .io_data_1_in_bits(PE_142_io_data_1_in_bits),
    .io_data_1_out_valid(PE_142_io_data_1_out_valid),
    .io_data_1_out_bits(PE_142_io_data_1_out_bits),
    .io_data_0_in_valid(PE_142_io_data_0_in_valid),
    .io_data_0_in_bits(PE_142_io_data_0_in_bits),
    .io_data_0_out_valid(PE_142_io_data_0_out_valid),
    .io_data_0_out_bits(PE_142_io_data_0_out_bits)
  );
  PE PE_143 ( // @[pe.scala 187:13]
    .clock(PE_143_clock),
    .reset(PE_143_reset),
    .io_data_2_out_valid(PE_143_io_data_2_out_valid),
    .io_data_2_out_bits(PE_143_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_143_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_143_io_data_1_in_valid),
    .io_data_1_in_bits(PE_143_io_data_1_in_bits),
    .io_data_1_out_valid(PE_143_io_data_1_out_valid),
    .io_data_1_out_bits(PE_143_io_data_1_out_bits),
    .io_data_0_in_valid(PE_143_io_data_0_in_valid),
    .io_data_0_in_bits(PE_143_io_data_0_in_bits),
    .io_data_0_out_valid(PE_143_io_data_0_out_valid),
    .io_data_0_out_bits(PE_143_io_data_0_out_bits)
  );
  PE PE_144 ( // @[pe.scala 187:13]
    .clock(PE_144_clock),
    .reset(PE_144_reset),
    .io_data_2_out_valid(PE_144_io_data_2_out_valid),
    .io_data_2_out_bits(PE_144_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_144_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_144_io_data_1_in_valid),
    .io_data_1_in_bits(PE_144_io_data_1_in_bits),
    .io_data_1_out_valid(PE_144_io_data_1_out_valid),
    .io_data_1_out_bits(PE_144_io_data_1_out_bits),
    .io_data_0_in_valid(PE_144_io_data_0_in_valid),
    .io_data_0_in_bits(PE_144_io_data_0_in_bits),
    .io_data_0_out_valid(PE_144_io_data_0_out_valid),
    .io_data_0_out_bits(PE_144_io_data_0_out_bits)
  );
  PE PE_145 ( // @[pe.scala 187:13]
    .clock(PE_145_clock),
    .reset(PE_145_reset),
    .io_data_2_out_valid(PE_145_io_data_2_out_valid),
    .io_data_2_out_bits(PE_145_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_145_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_145_io_data_1_in_valid),
    .io_data_1_in_bits(PE_145_io_data_1_in_bits),
    .io_data_1_out_valid(PE_145_io_data_1_out_valid),
    .io_data_1_out_bits(PE_145_io_data_1_out_bits),
    .io_data_0_in_valid(PE_145_io_data_0_in_valid),
    .io_data_0_in_bits(PE_145_io_data_0_in_bits),
    .io_data_0_out_valid(PE_145_io_data_0_out_valid),
    .io_data_0_out_bits(PE_145_io_data_0_out_bits)
  );
  PE PE_146 ( // @[pe.scala 187:13]
    .clock(PE_146_clock),
    .reset(PE_146_reset),
    .io_data_2_out_valid(PE_146_io_data_2_out_valid),
    .io_data_2_out_bits(PE_146_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_146_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_146_io_data_1_in_valid),
    .io_data_1_in_bits(PE_146_io_data_1_in_bits),
    .io_data_1_out_valid(PE_146_io_data_1_out_valid),
    .io_data_1_out_bits(PE_146_io_data_1_out_bits),
    .io_data_0_in_valid(PE_146_io_data_0_in_valid),
    .io_data_0_in_bits(PE_146_io_data_0_in_bits),
    .io_data_0_out_valid(PE_146_io_data_0_out_valid),
    .io_data_0_out_bits(PE_146_io_data_0_out_bits)
  );
  PE PE_147 ( // @[pe.scala 187:13]
    .clock(PE_147_clock),
    .reset(PE_147_reset),
    .io_data_2_out_valid(PE_147_io_data_2_out_valid),
    .io_data_2_out_bits(PE_147_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_147_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_147_io_data_1_in_valid),
    .io_data_1_in_bits(PE_147_io_data_1_in_bits),
    .io_data_1_out_valid(PE_147_io_data_1_out_valid),
    .io_data_1_out_bits(PE_147_io_data_1_out_bits),
    .io_data_0_in_valid(PE_147_io_data_0_in_valid),
    .io_data_0_in_bits(PE_147_io_data_0_in_bits),
    .io_data_0_out_valid(PE_147_io_data_0_out_valid),
    .io_data_0_out_bits(PE_147_io_data_0_out_bits)
  );
  PE PE_148 ( // @[pe.scala 187:13]
    .clock(PE_148_clock),
    .reset(PE_148_reset),
    .io_data_2_out_valid(PE_148_io_data_2_out_valid),
    .io_data_2_out_bits(PE_148_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_148_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_148_io_data_1_in_valid),
    .io_data_1_in_bits(PE_148_io_data_1_in_bits),
    .io_data_1_out_valid(PE_148_io_data_1_out_valid),
    .io_data_1_out_bits(PE_148_io_data_1_out_bits),
    .io_data_0_in_valid(PE_148_io_data_0_in_valid),
    .io_data_0_in_bits(PE_148_io_data_0_in_bits),
    .io_data_0_out_valid(PE_148_io_data_0_out_valid),
    .io_data_0_out_bits(PE_148_io_data_0_out_bits)
  );
  PE PE_149 ( // @[pe.scala 187:13]
    .clock(PE_149_clock),
    .reset(PE_149_reset),
    .io_data_2_out_valid(PE_149_io_data_2_out_valid),
    .io_data_2_out_bits(PE_149_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_149_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_149_io_data_1_in_valid),
    .io_data_1_in_bits(PE_149_io_data_1_in_bits),
    .io_data_1_out_valid(PE_149_io_data_1_out_valid),
    .io_data_1_out_bits(PE_149_io_data_1_out_bits),
    .io_data_0_in_valid(PE_149_io_data_0_in_valid),
    .io_data_0_in_bits(PE_149_io_data_0_in_bits),
    .io_data_0_out_valid(PE_149_io_data_0_out_valid),
    .io_data_0_out_bits(PE_149_io_data_0_out_bits)
  );
  PE PE_150 ( // @[pe.scala 187:13]
    .clock(PE_150_clock),
    .reset(PE_150_reset),
    .io_data_2_out_valid(PE_150_io_data_2_out_valid),
    .io_data_2_out_bits(PE_150_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_150_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_150_io_data_1_in_valid),
    .io_data_1_in_bits(PE_150_io_data_1_in_bits),
    .io_data_1_out_valid(PE_150_io_data_1_out_valid),
    .io_data_1_out_bits(PE_150_io_data_1_out_bits),
    .io_data_0_in_valid(PE_150_io_data_0_in_valid),
    .io_data_0_in_bits(PE_150_io_data_0_in_bits),
    .io_data_0_out_valid(PE_150_io_data_0_out_valid),
    .io_data_0_out_bits(PE_150_io_data_0_out_bits)
  );
  PE PE_151 ( // @[pe.scala 187:13]
    .clock(PE_151_clock),
    .reset(PE_151_reset),
    .io_data_2_out_valid(PE_151_io_data_2_out_valid),
    .io_data_2_out_bits(PE_151_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_151_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_151_io_data_1_in_valid),
    .io_data_1_in_bits(PE_151_io_data_1_in_bits),
    .io_data_1_out_valid(PE_151_io_data_1_out_valid),
    .io_data_1_out_bits(PE_151_io_data_1_out_bits),
    .io_data_0_in_valid(PE_151_io_data_0_in_valid),
    .io_data_0_in_bits(PE_151_io_data_0_in_bits),
    .io_data_0_out_valid(PE_151_io_data_0_out_valid),
    .io_data_0_out_bits(PE_151_io_data_0_out_bits)
  );
  PE PE_152 ( // @[pe.scala 187:13]
    .clock(PE_152_clock),
    .reset(PE_152_reset),
    .io_data_2_out_valid(PE_152_io_data_2_out_valid),
    .io_data_2_out_bits(PE_152_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_152_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_152_io_data_1_in_valid),
    .io_data_1_in_bits(PE_152_io_data_1_in_bits),
    .io_data_1_out_valid(PE_152_io_data_1_out_valid),
    .io_data_1_out_bits(PE_152_io_data_1_out_bits),
    .io_data_0_in_valid(PE_152_io_data_0_in_valid),
    .io_data_0_in_bits(PE_152_io_data_0_in_bits),
    .io_data_0_out_valid(PE_152_io_data_0_out_valid),
    .io_data_0_out_bits(PE_152_io_data_0_out_bits)
  );
  PE PE_153 ( // @[pe.scala 187:13]
    .clock(PE_153_clock),
    .reset(PE_153_reset),
    .io_data_2_out_valid(PE_153_io_data_2_out_valid),
    .io_data_2_out_bits(PE_153_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_153_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_153_io_data_1_in_valid),
    .io_data_1_in_bits(PE_153_io_data_1_in_bits),
    .io_data_1_out_valid(PE_153_io_data_1_out_valid),
    .io_data_1_out_bits(PE_153_io_data_1_out_bits),
    .io_data_0_in_valid(PE_153_io_data_0_in_valid),
    .io_data_0_in_bits(PE_153_io_data_0_in_bits),
    .io_data_0_out_valid(PE_153_io_data_0_out_valid),
    .io_data_0_out_bits(PE_153_io_data_0_out_bits)
  );
  PE PE_154 ( // @[pe.scala 187:13]
    .clock(PE_154_clock),
    .reset(PE_154_reset),
    .io_data_2_out_valid(PE_154_io_data_2_out_valid),
    .io_data_2_out_bits(PE_154_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_154_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_154_io_data_1_in_valid),
    .io_data_1_in_bits(PE_154_io_data_1_in_bits),
    .io_data_1_out_valid(PE_154_io_data_1_out_valid),
    .io_data_1_out_bits(PE_154_io_data_1_out_bits),
    .io_data_0_in_valid(PE_154_io_data_0_in_valid),
    .io_data_0_in_bits(PE_154_io_data_0_in_bits),
    .io_data_0_out_valid(PE_154_io_data_0_out_valid),
    .io_data_0_out_bits(PE_154_io_data_0_out_bits)
  );
  PE PE_155 ( // @[pe.scala 187:13]
    .clock(PE_155_clock),
    .reset(PE_155_reset),
    .io_data_2_out_valid(PE_155_io_data_2_out_valid),
    .io_data_2_out_bits(PE_155_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_155_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_155_io_data_1_in_valid),
    .io_data_1_in_bits(PE_155_io_data_1_in_bits),
    .io_data_1_out_valid(PE_155_io_data_1_out_valid),
    .io_data_1_out_bits(PE_155_io_data_1_out_bits),
    .io_data_0_in_valid(PE_155_io_data_0_in_valid),
    .io_data_0_in_bits(PE_155_io_data_0_in_bits),
    .io_data_0_out_valid(PE_155_io_data_0_out_valid),
    .io_data_0_out_bits(PE_155_io_data_0_out_bits)
  );
  PE PE_156 ( // @[pe.scala 187:13]
    .clock(PE_156_clock),
    .reset(PE_156_reset),
    .io_data_2_out_valid(PE_156_io_data_2_out_valid),
    .io_data_2_out_bits(PE_156_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_156_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_156_io_data_1_in_valid),
    .io_data_1_in_bits(PE_156_io_data_1_in_bits),
    .io_data_1_out_valid(PE_156_io_data_1_out_valid),
    .io_data_1_out_bits(PE_156_io_data_1_out_bits),
    .io_data_0_in_valid(PE_156_io_data_0_in_valid),
    .io_data_0_in_bits(PE_156_io_data_0_in_bits),
    .io_data_0_out_valid(PE_156_io_data_0_out_valid),
    .io_data_0_out_bits(PE_156_io_data_0_out_bits)
  );
  PE PE_157 ( // @[pe.scala 187:13]
    .clock(PE_157_clock),
    .reset(PE_157_reset),
    .io_data_2_out_valid(PE_157_io_data_2_out_valid),
    .io_data_2_out_bits(PE_157_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_157_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_157_io_data_1_in_valid),
    .io_data_1_in_bits(PE_157_io_data_1_in_bits),
    .io_data_1_out_valid(PE_157_io_data_1_out_valid),
    .io_data_1_out_bits(PE_157_io_data_1_out_bits),
    .io_data_0_in_valid(PE_157_io_data_0_in_valid),
    .io_data_0_in_bits(PE_157_io_data_0_in_bits),
    .io_data_0_out_valid(PE_157_io_data_0_out_valid),
    .io_data_0_out_bits(PE_157_io_data_0_out_bits)
  );
  PE PE_158 ( // @[pe.scala 187:13]
    .clock(PE_158_clock),
    .reset(PE_158_reset),
    .io_data_2_out_valid(PE_158_io_data_2_out_valid),
    .io_data_2_out_bits(PE_158_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_158_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_158_io_data_1_in_valid),
    .io_data_1_in_bits(PE_158_io_data_1_in_bits),
    .io_data_1_out_valid(PE_158_io_data_1_out_valid),
    .io_data_1_out_bits(PE_158_io_data_1_out_bits),
    .io_data_0_in_valid(PE_158_io_data_0_in_valid),
    .io_data_0_in_bits(PE_158_io_data_0_in_bits),
    .io_data_0_out_valid(PE_158_io_data_0_out_valid),
    .io_data_0_out_bits(PE_158_io_data_0_out_bits)
  );
  PE PE_159 ( // @[pe.scala 187:13]
    .clock(PE_159_clock),
    .reset(PE_159_reset),
    .io_data_2_out_valid(PE_159_io_data_2_out_valid),
    .io_data_2_out_bits(PE_159_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_159_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_159_io_data_1_in_valid),
    .io_data_1_in_bits(PE_159_io_data_1_in_bits),
    .io_data_1_out_valid(PE_159_io_data_1_out_valid),
    .io_data_1_out_bits(PE_159_io_data_1_out_bits),
    .io_data_0_in_valid(PE_159_io_data_0_in_valid),
    .io_data_0_in_bits(PE_159_io_data_0_in_bits),
    .io_data_0_out_valid(PE_159_io_data_0_out_valid),
    .io_data_0_out_bits(PE_159_io_data_0_out_bits)
  );
  PE PE_160 ( // @[pe.scala 187:13]
    .clock(PE_160_clock),
    .reset(PE_160_reset),
    .io_data_2_out_valid(PE_160_io_data_2_out_valid),
    .io_data_2_out_bits(PE_160_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_160_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_160_io_data_1_in_valid),
    .io_data_1_in_bits(PE_160_io_data_1_in_bits),
    .io_data_1_out_valid(PE_160_io_data_1_out_valid),
    .io_data_1_out_bits(PE_160_io_data_1_out_bits),
    .io_data_0_in_valid(PE_160_io_data_0_in_valid),
    .io_data_0_in_bits(PE_160_io_data_0_in_bits),
    .io_data_0_out_valid(PE_160_io_data_0_out_valid),
    .io_data_0_out_bits(PE_160_io_data_0_out_bits)
  );
  PE PE_161 ( // @[pe.scala 187:13]
    .clock(PE_161_clock),
    .reset(PE_161_reset),
    .io_data_2_out_valid(PE_161_io_data_2_out_valid),
    .io_data_2_out_bits(PE_161_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_161_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_161_io_data_1_in_valid),
    .io_data_1_in_bits(PE_161_io_data_1_in_bits),
    .io_data_1_out_valid(PE_161_io_data_1_out_valid),
    .io_data_1_out_bits(PE_161_io_data_1_out_bits),
    .io_data_0_in_valid(PE_161_io_data_0_in_valid),
    .io_data_0_in_bits(PE_161_io_data_0_in_bits),
    .io_data_0_out_valid(PE_161_io_data_0_out_valid),
    .io_data_0_out_bits(PE_161_io_data_0_out_bits)
  );
  PE PE_162 ( // @[pe.scala 187:13]
    .clock(PE_162_clock),
    .reset(PE_162_reset),
    .io_data_2_out_valid(PE_162_io_data_2_out_valid),
    .io_data_2_out_bits(PE_162_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_162_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_162_io_data_1_in_valid),
    .io_data_1_in_bits(PE_162_io_data_1_in_bits),
    .io_data_1_out_valid(PE_162_io_data_1_out_valid),
    .io_data_1_out_bits(PE_162_io_data_1_out_bits),
    .io_data_0_in_valid(PE_162_io_data_0_in_valid),
    .io_data_0_in_bits(PE_162_io_data_0_in_bits),
    .io_data_0_out_valid(PE_162_io_data_0_out_valid),
    .io_data_0_out_bits(PE_162_io_data_0_out_bits)
  );
  PE PE_163 ( // @[pe.scala 187:13]
    .clock(PE_163_clock),
    .reset(PE_163_reset),
    .io_data_2_out_valid(PE_163_io_data_2_out_valid),
    .io_data_2_out_bits(PE_163_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_163_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_163_io_data_1_in_valid),
    .io_data_1_in_bits(PE_163_io_data_1_in_bits),
    .io_data_1_out_valid(PE_163_io_data_1_out_valid),
    .io_data_1_out_bits(PE_163_io_data_1_out_bits),
    .io_data_0_in_valid(PE_163_io_data_0_in_valid),
    .io_data_0_in_bits(PE_163_io_data_0_in_bits),
    .io_data_0_out_valid(PE_163_io_data_0_out_valid),
    .io_data_0_out_bits(PE_163_io_data_0_out_bits)
  );
  PE PE_164 ( // @[pe.scala 187:13]
    .clock(PE_164_clock),
    .reset(PE_164_reset),
    .io_data_2_out_valid(PE_164_io_data_2_out_valid),
    .io_data_2_out_bits(PE_164_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_164_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_164_io_data_1_in_valid),
    .io_data_1_in_bits(PE_164_io_data_1_in_bits),
    .io_data_1_out_valid(PE_164_io_data_1_out_valid),
    .io_data_1_out_bits(PE_164_io_data_1_out_bits),
    .io_data_0_in_valid(PE_164_io_data_0_in_valid),
    .io_data_0_in_bits(PE_164_io_data_0_in_bits),
    .io_data_0_out_valid(PE_164_io_data_0_out_valid),
    .io_data_0_out_bits(PE_164_io_data_0_out_bits)
  );
  PE PE_165 ( // @[pe.scala 187:13]
    .clock(PE_165_clock),
    .reset(PE_165_reset),
    .io_data_2_out_valid(PE_165_io_data_2_out_valid),
    .io_data_2_out_bits(PE_165_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_165_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_165_io_data_1_in_valid),
    .io_data_1_in_bits(PE_165_io_data_1_in_bits),
    .io_data_1_out_valid(PE_165_io_data_1_out_valid),
    .io_data_1_out_bits(PE_165_io_data_1_out_bits),
    .io_data_0_in_valid(PE_165_io_data_0_in_valid),
    .io_data_0_in_bits(PE_165_io_data_0_in_bits),
    .io_data_0_out_valid(PE_165_io_data_0_out_valid),
    .io_data_0_out_bits(PE_165_io_data_0_out_bits)
  );
  PE PE_166 ( // @[pe.scala 187:13]
    .clock(PE_166_clock),
    .reset(PE_166_reset),
    .io_data_2_out_valid(PE_166_io_data_2_out_valid),
    .io_data_2_out_bits(PE_166_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_166_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_166_io_data_1_in_valid),
    .io_data_1_in_bits(PE_166_io_data_1_in_bits),
    .io_data_1_out_valid(PE_166_io_data_1_out_valid),
    .io_data_1_out_bits(PE_166_io_data_1_out_bits),
    .io_data_0_in_valid(PE_166_io_data_0_in_valid),
    .io_data_0_in_bits(PE_166_io_data_0_in_bits),
    .io_data_0_out_valid(PE_166_io_data_0_out_valid),
    .io_data_0_out_bits(PE_166_io_data_0_out_bits)
  );
  PE PE_167 ( // @[pe.scala 187:13]
    .clock(PE_167_clock),
    .reset(PE_167_reset),
    .io_data_2_out_valid(PE_167_io_data_2_out_valid),
    .io_data_2_out_bits(PE_167_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_167_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_167_io_data_1_in_valid),
    .io_data_1_in_bits(PE_167_io_data_1_in_bits),
    .io_data_1_out_valid(PE_167_io_data_1_out_valid),
    .io_data_1_out_bits(PE_167_io_data_1_out_bits),
    .io_data_0_in_valid(PE_167_io_data_0_in_valid),
    .io_data_0_in_bits(PE_167_io_data_0_in_bits),
    .io_data_0_out_valid(PE_167_io_data_0_out_valid),
    .io_data_0_out_bits(PE_167_io_data_0_out_bits)
  );
  PE PE_168 ( // @[pe.scala 187:13]
    .clock(PE_168_clock),
    .reset(PE_168_reset),
    .io_data_2_out_valid(PE_168_io_data_2_out_valid),
    .io_data_2_out_bits(PE_168_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_168_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_168_io_data_1_in_valid),
    .io_data_1_in_bits(PE_168_io_data_1_in_bits),
    .io_data_1_out_valid(PE_168_io_data_1_out_valid),
    .io_data_1_out_bits(PE_168_io_data_1_out_bits),
    .io_data_0_in_valid(PE_168_io_data_0_in_valid),
    .io_data_0_in_bits(PE_168_io_data_0_in_bits),
    .io_data_0_out_valid(PE_168_io_data_0_out_valid),
    .io_data_0_out_bits(PE_168_io_data_0_out_bits)
  );
  PE PE_169 ( // @[pe.scala 187:13]
    .clock(PE_169_clock),
    .reset(PE_169_reset),
    .io_data_2_out_valid(PE_169_io_data_2_out_valid),
    .io_data_2_out_bits(PE_169_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_169_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_169_io_data_1_in_valid),
    .io_data_1_in_bits(PE_169_io_data_1_in_bits),
    .io_data_1_out_valid(PE_169_io_data_1_out_valid),
    .io_data_1_out_bits(PE_169_io_data_1_out_bits),
    .io_data_0_in_valid(PE_169_io_data_0_in_valid),
    .io_data_0_in_bits(PE_169_io_data_0_in_bits),
    .io_data_0_out_valid(PE_169_io_data_0_out_valid),
    .io_data_0_out_bits(PE_169_io_data_0_out_bits)
  );
  PE PE_170 ( // @[pe.scala 187:13]
    .clock(PE_170_clock),
    .reset(PE_170_reset),
    .io_data_2_out_valid(PE_170_io_data_2_out_valid),
    .io_data_2_out_bits(PE_170_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_170_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_170_io_data_1_in_valid),
    .io_data_1_in_bits(PE_170_io_data_1_in_bits),
    .io_data_1_out_valid(PE_170_io_data_1_out_valid),
    .io_data_1_out_bits(PE_170_io_data_1_out_bits),
    .io_data_0_in_valid(PE_170_io_data_0_in_valid),
    .io_data_0_in_bits(PE_170_io_data_0_in_bits),
    .io_data_0_out_valid(PE_170_io_data_0_out_valid),
    .io_data_0_out_bits(PE_170_io_data_0_out_bits)
  );
  PE PE_171 ( // @[pe.scala 187:13]
    .clock(PE_171_clock),
    .reset(PE_171_reset),
    .io_data_2_out_valid(PE_171_io_data_2_out_valid),
    .io_data_2_out_bits(PE_171_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_171_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_171_io_data_1_in_valid),
    .io_data_1_in_bits(PE_171_io_data_1_in_bits),
    .io_data_1_out_valid(PE_171_io_data_1_out_valid),
    .io_data_1_out_bits(PE_171_io_data_1_out_bits),
    .io_data_0_in_valid(PE_171_io_data_0_in_valid),
    .io_data_0_in_bits(PE_171_io_data_0_in_bits),
    .io_data_0_out_valid(PE_171_io_data_0_out_valid),
    .io_data_0_out_bits(PE_171_io_data_0_out_bits)
  );
  PE PE_172 ( // @[pe.scala 187:13]
    .clock(PE_172_clock),
    .reset(PE_172_reset),
    .io_data_2_out_valid(PE_172_io_data_2_out_valid),
    .io_data_2_out_bits(PE_172_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_172_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_172_io_data_1_in_valid),
    .io_data_1_in_bits(PE_172_io_data_1_in_bits),
    .io_data_1_out_valid(PE_172_io_data_1_out_valid),
    .io_data_1_out_bits(PE_172_io_data_1_out_bits),
    .io_data_0_in_valid(PE_172_io_data_0_in_valid),
    .io_data_0_in_bits(PE_172_io_data_0_in_bits),
    .io_data_0_out_valid(PE_172_io_data_0_out_valid),
    .io_data_0_out_bits(PE_172_io_data_0_out_bits)
  );
  PE PE_173 ( // @[pe.scala 187:13]
    .clock(PE_173_clock),
    .reset(PE_173_reset),
    .io_data_2_out_valid(PE_173_io_data_2_out_valid),
    .io_data_2_out_bits(PE_173_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_173_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_173_io_data_1_in_valid),
    .io_data_1_in_bits(PE_173_io_data_1_in_bits),
    .io_data_1_out_valid(PE_173_io_data_1_out_valid),
    .io_data_1_out_bits(PE_173_io_data_1_out_bits),
    .io_data_0_in_valid(PE_173_io_data_0_in_valid),
    .io_data_0_in_bits(PE_173_io_data_0_in_bits),
    .io_data_0_out_valid(PE_173_io_data_0_out_valid),
    .io_data_0_out_bits(PE_173_io_data_0_out_bits)
  );
  PE PE_174 ( // @[pe.scala 187:13]
    .clock(PE_174_clock),
    .reset(PE_174_reset),
    .io_data_2_out_valid(PE_174_io_data_2_out_valid),
    .io_data_2_out_bits(PE_174_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_174_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_174_io_data_1_in_valid),
    .io_data_1_in_bits(PE_174_io_data_1_in_bits),
    .io_data_1_out_valid(PE_174_io_data_1_out_valid),
    .io_data_1_out_bits(PE_174_io_data_1_out_bits),
    .io_data_0_in_valid(PE_174_io_data_0_in_valid),
    .io_data_0_in_bits(PE_174_io_data_0_in_bits),
    .io_data_0_out_valid(PE_174_io_data_0_out_valid),
    .io_data_0_out_bits(PE_174_io_data_0_out_bits)
  );
  PE PE_175 ( // @[pe.scala 187:13]
    .clock(PE_175_clock),
    .reset(PE_175_reset),
    .io_data_2_out_valid(PE_175_io_data_2_out_valid),
    .io_data_2_out_bits(PE_175_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_175_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_175_io_data_1_in_valid),
    .io_data_1_in_bits(PE_175_io_data_1_in_bits),
    .io_data_1_out_valid(PE_175_io_data_1_out_valid),
    .io_data_1_out_bits(PE_175_io_data_1_out_bits),
    .io_data_0_in_valid(PE_175_io_data_0_in_valid),
    .io_data_0_in_bits(PE_175_io_data_0_in_bits),
    .io_data_0_out_valid(PE_175_io_data_0_out_valid),
    .io_data_0_out_bits(PE_175_io_data_0_out_bits)
  );
  PE PE_176 ( // @[pe.scala 187:13]
    .clock(PE_176_clock),
    .reset(PE_176_reset),
    .io_data_2_out_valid(PE_176_io_data_2_out_valid),
    .io_data_2_out_bits(PE_176_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_176_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_176_io_data_1_in_valid),
    .io_data_1_in_bits(PE_176_io_data_1_in_bits),
    .io_data_1_out_valid(PE_176_io_data_1_out_valid),
    .io_data_1_out_bits(PE_176_io_data_1_out_bits),
    .io_data_0_in_valid(PE_176_io_data_0_in_valid),
    .io_data_0_in_bits(PE_176_io_data_0_in_bits),
    .io_data_0_out_valid(PE_176_io_data_0_out_valid),
    .io_data_0_out_bits(PE_176_io_data_0_out_bits)
  );
  PE PE_177 ( // @[pe.scala 187:13]
    .clock(PE_177_clock),
    .reset(PE_177_reset),
    .io_data_2_out_valid(PE_177_io_data_2_out_valid),
    .io_data_2_out_bits(PE_177_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_177_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_177_io_data_1_in_valid),
    .io_data_1_in_bits(PE_177_io_data_1_in_bits),
    .io_data_1_out_valid(PE_177_io_data_1_out_valid),
    .io_data_1_out_bits(PE_177_io_data_1_out_bits),
    .io_data_0_in_valid(PE_177_io_data_0_in_valid),
    .io_data_0_in_bits(PE_177_io_data_0_in_bits),
    .io_data_0_out_valid(PE_177_io_data_0_out_valid),
    .io_data_0_out_bits(PE_177_io_data_0_out_bits)
  );
  PE PE_178 ( // @[pe.scala 187:13]
    .clock(PE_178_clock),
    .reset(PE_178_reset),
    .io_data_2_out_valid(PE_178_io_data_2_out_valid),
    .io_data_2_out_bits(PE_178_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_178_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_178_io_data_1_in_valid),
    .io_data_1_in_bits(PE_178_io_data_1_in_bits),
    .io_data_1_out_valid(PE_178_io_data_1_out_valid),
    .io_data_1_out_bits(PE_178_io_data_1_out_bits),
    .io_data_0_in_valid(PE_178_io_data_0_in_valid),
    .io_data_0_in_bits(PE_178_io_data_0_in_bits),
    .io_data_0_out_valid(PE_178_io_data_0_out_valid),
    .io_data_0_out_bits(PE_178_io_data_0_out_bits)
  );
  PE PE_179 ( // @[pe.scala 187:13]
    .clock(PE_179_clock),
    .reset(PE_179_reset),
    .io_data_2_out_valid(PE_179_io_data_2_out_valid),
    .io_data_2_out_bits(PE_179_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_179_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_179_io_data_1_in_valid),
    .io_data_1_in_bits(PE_179_io_data_1_in_bits),
    .io_data_1_out_valid(PE_179_io_data_1_out_valid),
    .io_data_1_out_bits(PE_179_io_data_1_out_bits),
    .io_data_0_in_valid(PE_179_io_data_0_in_valid),
    .io_data_0_in_bits(PE_179_io_data_0_in_bits),
    .io_data_0_out_valid(PE_179_io_data_0_out_valid),
    .io_data_0_out_bits(PE_179_io_data_0_out_bits)
  );
  PE PE_180 ( // @[pe.scala 187:13]
    .clock(PE_180_clock),
    .reset(PE_180_reset),
    .io_data_2_out_valid(PE_180_io_data_2_out_valid),
    .io_data_2_out_bits(PE_180_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_180_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_180_io_data_1_in_valid),
    .io_data_1_in_bits(PE_180_io_data_1_in_bits),
    .io_data_1_out_valid(PE_180_io_data_1_out_valid),
    .io_data_1_out_bits(PE_180_io_data_1_out_bits),
    .io_data_0_in_valid(PE_180_io_data_0_in_valid),
    .io_data_0_in_bits(PE_180_io_data_0_in_bits),
    .io_data_0_out_valid(PE_180_io_data_0_out_valid),
    .io_data_0_out_bits(PE_180_io_data_0_out_bits)
  );
  PE PE_181 ( // @[pe.scala 187:13]
    .clock(PE_181_clock),
    .reset(PE_181_reset),
    .io_data_2_out_valid(PE_181_io_data_2_out_valid),
    .io_data_2_out_bits(PE_181_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_181_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_181_io_data_1_in_valid),
    .io_data_1_in_bits(PE_181_io_data_1_in_bits),
    .io_data_1_out_valid(PE_181_io_data_1_out_valid),
    .io_data_1_out_bits(PE_181_io_data_1_out_bits),
    .io_data_0_in_valid(PE_181_io_data_0_in_valid),
    .io_data_0_in_bits(PE_181_io_data_0_in_bits),
    .io_data_0_out_valid(PE_181_io_data_0_out_valid),
    .io_data_0_out_bits(PE_181_io_data_0_out_bits)
  );
  PE PE_182 ( // @[pe.scala 187:13]
    .clock(PE_182_clock),
    .reset(PE_182_reset),
    .io_data_2_out_valid(PE_182_io_data_2_out_valid),
    .io_data_2_out_bits(PE_182_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_182_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_182_io_data_1_in_valid),
    .io_data_1_in_bits(PE_182_io_data_1_in_bits),
    .io_data_1_out_valid(PE_182_io_data_1_out_valid),
    .io_data_1_out_bits(PE_182_io_data_1_out_bits),
    .io_data_0_in_valid(PE_182_io_data_0_in_valid),
    .io_data_0_in_bits(PE_182_io_data_0_in_bits),
    .io_data_0_out_valid(PE_182_io_data_0_out_valid),
    .io_data_0_out_bits(PE_182_io_data_0_out_bits)
  );
  PE PE_183 ( // @[pe.scala 187:13]
    .clock(PE_183_clock),
    .reset(PE_183_reset),
    .io_data_2_out_valid(PE_183_io_data_2_out_valid),
    .io_data_2_out_bits(PE_183_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_183_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_183_io_data_1_in_valid),
    .io_data_1_in_bits(PE_183_io_data_1_in_bits),
    .io_data_1_out_valid(PE_183_io_data_1_out_valid),
    .io_data_1_out_bits(PE_183_io_data_1_out_bits),
    .io_data_0_in_valid(PE_183_io_data_0_in_valid),
    .io_data_0_in_bits(PE_183_io_data_0_in_bits),
    .io_data_0_out_valid(PE_183_io_data_0_out_valid),
    .io_data_0_out_bits(PE_183_io_data_0_out_bits)
  );
  PE PE_184 ( // @[pe.scala 187:13]
    .clock(PE_184_clock),
    .reset(PE_184_reset),
    .io_data_2_out_valid(PE_184_io_data_2_out_valid),
    .io_data_2_out_bits(PE_184_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_184_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_184_io_data_1_in_valid),
    .io_data_1_in_bits(PE_184_io_data_1_in_bits),
    .io_data_1_out_valid(PE_184_io_data_1_out_valid),
    .io_data_1_out_bits(PE_184_io_data_1_out_bits),
    .io_data_0_in_valid(PE_184_io_data_0_in_valid),
    .io_data_0_in_bits(PE_184_io_data_0_in_bits),
    .io_data_0_out_valid(PE_184_io_data_0_out_valid),
    .io_data_0_out_bits(PE_184_io_data_0_out_bits)
  );
  PE PE_185 ( // @[pe.scala 187:13]
    .clock(PE_185_clock),
    .reset(PE_185_reset),
    .io_data_2_out_valid(PE_185_io_data_2_out_valid),
    .io_data_2_out_bits(PE_185_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_185_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_185_io_data_1_in_valid),
    .io_data_1_in_bits(PE_185_io_data_1_in_bits),
    .io_data_1_out_valid(PE_185_io_data_1_out_valid),
    .io_data_1_out_bits(PE_185_io_data_1_out_bits),
    .io_data_0_in_valid(PE_185_io_data_0_in_valid),
    .io_data_0_in_bits(PE_185_io_data_0_in_bits),
    .io_data_0_out_valid(PE_185_io_data_0_out_valid),
    .io_data_0_out_bits(PE_185_io_data_0_out_bits)
  );
  PE PE_186 ( // @[pe.scala 187:13]
    .clock(PE_186_clock),
    .reset(PE_186_reset),
    .io_data_2_out_valid(PE_186_io_data_2_out_valid),
    .io_data_2_out_bits(PE_186_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_186_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_186_io_data_1_in_valid),
    .io_data_1_in_bits(PE_186_io_data_1_in_bits),
    .io_data_1_out_valid(PE_186_io_data_1_out_valid),
    .io_data_1_out_bits(PE_186_io_data_1_out_bits),
    .io_data_0_in_valid(PE_186_io_data_0_in_valid),
    .io_data_0_in_bits(PE_186_io_data_0_in_bits),
    .io_data_0_out_valid(PE_186_io_data_0_out_valid),
    .io_data_0_out_bits(PE_186_io_data_0_out_bits)
  );
  PE PE_187 ( // @[pe.scala 187:13]
    .clock(PE_187_clock),
    .reset(PE_187_reset),
    .io_data_2_out_valid(PE_187_io_data_2_out_valid),
    .io_data_2_out_bits(PE_187_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_187_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_187_io_data_1_in_valid),
    .io_data_1_in_bits(PE_187_io_data_1_in_bits),
    .io_data_1_out_valid(PE_187_io_data_1_out_valid),
    .io_data_1_out_bits(PE_187_io_data_1_out_bits),
    .io_data_0_in_valid(PE_187_io_data_0_in_valid),
    .io_data_0_in_bits(PE_187_io_data_0_in_bits),
    .io_data_0_out_valid(PE_187_io_data_0_out_valid),
    .io_data_0_out_bits(PE_187_io_data_0_out_bits)
  );
  PE PE_188 ( // @[pe.scala 187:13]
    .clock(PE_188_clock),
    .reset(PE_188_reset),
    .io_data_2_out_valid(PE_188_io_data_2_out_valid),
    .io_data_2_out_bits(PE_188_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_188_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_188_io_data_1_in_valid),
    .io_data_1_in_bits(PE_188_io_data_1_in_bits),
    .io_data_1_out_valid(PE_188_io_data_1_out_valid),
    .io_data_1_out_bits(PE_188_io_data_1_out_bits),
    .io_data_0_in_valid(PE_188_io_data_0_in_valid),
    .io_data_0_in_bits(PE_188_io_data_0_in_bits),
    .io_data_0_out_valid(PE_188_io_data_0_out_valid),
    .io_data_0_out_bits(PE_188_io_data_0_out_bits)
  );
  PE PE_189 ( // @[pe.scala 187:13]
    .clock(PE_189_clock),
    .reset(PE_189_reset),
    .io_data_2_out_valid(PE_189_io_data_2_out_valid),
    .io_data_2_out_bits(PE_189_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_189_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_189_io_data_1_in_valid),
    .io_data_1_in_bits(PE_189_io_data_1_in_bits),
    .io_data_1_out_valid(PE_189_io_data_1_out_valid),
    .io_data_1_out_bits(PE_189_io_data_1_out_bits),
    .io_data_0_in_valid(PE_189_io_data_0_in_valid),
    .io_data_0_in_bits(PE_189_io_data_0_in_bits),
    .io_data_0_out_valid(PE_189_io_data_0_out_valid),
    .io_data_0_out_bits(PE_189_io_data_0_out_bits)
  );
  PE PE_190 ( // @[pe.scala 187:13]
    .clock(PE_190_clock),
    .reset(PE_190_reset),
    .io_data_2_out_valid(PE_190_io_data_2_out_valid),
    .io_data_2_out_bits(PE_190_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_190_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_190_io_data_1_in_valid),
    .io_data_1_in_bits(PE_190_io_data_1_in_bits),
    .io_data_1_out_valid(PE_190_io_data_1_out_valid),
    .io_data_1_out_bits(PE_190_io_data_1_out_bits),
    .io_data_0_in_valid(PE_190_io_data_0_in_valid),
    .io_data_0_in_bits(PE_190_io_data_0_in_bits),
    .io_data_0_out_valid(PE_190_io_data_0_out_valid),
    .io_data_0_out_bits(PE_190_io_data_0_out_bits)
  );
  PE PE_191 ( // @[pe.scala 187:13]
    .clock(PE_191_clock),
    .reset(PE_191_reset),
    .io_data_2_out_valid(PE_191_io_data_2_out_valid),
    .io_data_2_out_bits(PE_191_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_191_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_191_io_data_1_in_valid),
    .io_data_1_in_bits(PE_191_io_data_1_in_bits),
    .io_data_1_out_valid(PE_191_io_data_1_out_valid),
    .io_data_1_out_bits(PE_191_io_data_1_out_bits),
    .io_data_0_in_valid(PE_191_io_data_0_in_valid),
    .io_data_0_in_bits(PE_191_io_data_0_in_bits),
    .io_data_0_out_valid(PE_191_io_data_0_out_valid),
    .io_data_0_out_bits(PE_191_io_data_0_out_bits)
  );
  PE PE_192 ( // @[pe.scala 187:13]
    .clock(PE_192_clock),
    .reset(PE_192_reset),
    .io_data_2_out_valid(PE_192_io_data_2_out_valid),
    .io_data_2_out_bits(PE_192_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_192_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_192_io_data_1_in_valid),
    .io_data_1_in_bits(PE_192_io_data_1_in_bits),
    .io_data_1_out_valid(PE_192_io_data_1_out_valid),
    .io_data_1_out_bits(PE_192_io_data_1_out_bits),
    .io_data_0_in_valid(PE_192_io_data_0_in_valid),
    .io_data_0_in_bits(PE_192_io_data_0_in_bits),
    .io_data_0_out_valid(PE_192_io_data_0_out_valid),
    .io_data_0_out_bits(PE_192_io_data_0_out_bits)
  );
  PE PE_193 ( // @[pe.scala 187:13]
    .clock(PE_193_clock),
    .reset(PE_193_reset),
    .io_data_2_out_valid(PE_193_io_data_2_out_valid),
    .io_data_2_out_bits(PE_193_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_193_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_193_io_data_1_in_valid),
    .io_data_1_in_bits(PE_193_io_data_1_in_bits),
    .io_data_1_out_valid(PE_193_io_data_1_out_valid),
    .io_data_1_out_bits(PE_193_io_data_1_out_bits),
    .io_data_0_in_valid(PE_193_io_data_0_in_valid),
    .io_data_0_in_bits(PE_193_io_data_0_in_bits),
    .io_data_0_out_valid(PE_193_io_data_0_out_valid),
    .io_data_0_out_bits(PE_193_io_data_0_out_bits)
  );
  PE PE_194 ( // @[pe.scala 187:13]
    .clock(PE_194_clock),
    .reset(PE_194_reset),
    .io_data_2_out_valid(PE_194_io_data_2_out_valid),
    .io_data_2_out_bits(PE_194_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_194_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_194_io_data_1_in_valid),
    .io_data_1_in_bits(PE_194_io_data_1_in_bits),
    .io_data_1_out_valid(PE_194_io_data_1_out_valid),
    .io_data_1_out_bits(PE_194_io_data_1_out_bits),
    .io_data_0_in_valid(PE_194_io_data_0_in_valid),
    .io_data_0_in_bits(PE_194_io_data_0_in_bits),
    .io_data_0_out_valid(PE_194_io_data_0_out_valid),
    .io_data_0_out_bits(PE_194_io_data_0_out_bits)
  );
  PE PE_195 ( // @[pe.scala 187:13]
    .clock(PE_195_clock),
    .reset(PE_195_reset),
    .io_data_2_out_valid(PE_195_io_data_2_out_valid),
    .io_data_2_out_bits(PE_195_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_195_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_195_io_data_1_in_valid),
    .io_data_1_in_bits(PE_195_io_data_1_in_bits),
    .io_data_1_out_valid(PE_195_io_data_1_out_valid),
    .io_data_1_out_bits(PE_195_io_data_1_out_bits),
    .io_data_0_in_valid(PE_195_io_data_0_in_valid),
    .io_data_0_in_bits(PE_195_io_data_0_in_bits),
    .io_data_0_out_valid(PE_195_io_data_0_out_valid),
    .io_data_0_out_bits(PE_195_io_data_0_out_bits)
  );
  PE PE_196 ( // @[pe.scala 187:13]
    .clock(PE_196_clock),
    .reset(PE_196_reset),
    .io_data_2_out_valid(PE_196_io_data_2_out_valid),
    .io_data_2_out_bits(PE_196_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_196_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_196_io_data_1_in_valid),
    .io_data_1_in_bits(PE_196_io_data_1_in_bits),
    .io_data_1_out_valid(PE_196_io_data_1_out_valid),
    .io_data_1_out_bits(PE_196_io_data_1_out_bits),
    .io_data_0_in_valid(PE_196_io_data_0_in_valid),
    .io_data_0_in_bits(PE_196_io_data_0_in_bits),
    .io_data_0_out_valid(PE_196_io_data_0_out_valid),
    .io_data_0_out_bits(PE_196_io_data_0_out_bits)
  );
  PE PE_197 ( // @[pe.scala 187:13]
    .clock(PE_197_clock),
    .reset(PE_197_reset),
    .io_data_2_out_valid(PE_197_io_data_2_out_valid),
    .io_data_2_out_bits(PE_197_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_197_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_197_io_data_1_in_valid),
    .io_data_1_in_bits(PE_197_io_data_1_in_bits),
    .io_data_1_out_valid(PE_197_io_data_1_out_valid),
    .io_data_1_out_bits(PE_197_io_data_1_out_bits),
    .io_data_0_in_valid(PE_197_io_data_0_in_valid),
    .io_data_0_in_bits(PE_197_io_data_0_in_bits),
    .io_data_0_out_valid(PE_197_io_data_0_out_valid),
    .io_data_0_out_bits(PE_197_io_data_0_out_bits)
  );
  PE PE_198 ( // @[pe.scala 187:13]
    .clock(PE_198_clock),
    .reset(PE_198_reset),
    .io_data_2_out_valid(PE_198_io_data_2_out_valid),
    .io_data_2_out_bits(PE_198_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_198_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_198_io_data_1_in_valid),
    .io_data_1_in_bits(PE_198_io_data_1_in_bits),
    .io_data_1_out_valid(PE_198_io_data_1_out_valid),
    .io_data_1_out_bits(PE_198_io_data_1_out_bits),
    .io_data_0_in_valid(PE_198_io_data_0_in_valid),
    .io_data_0_in_bits(PE_198_io_data_0_in_bits),
    .io_data_0_out_valid(PE_198_io_data_0_out_valid),
    .io_data_0_out_bits(PE_198_io_data_0_out_bits)
  );
  PE PE_199 ( // @[pe.scala 187:13]
    .clock(PE_199_clock),
    .reset(PE_199_reset),
    .io_data_2_out_valid(PE_199_io_data_2_out_valid),
    .io_data_2_out_bits(PE_199_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_199_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_199_io_data_1_in_valid),
    .io_data_1_in_bits(PE_199_io_data_1_in_bits),
    .io_data_1_out_valid(PE_199_io_data_1_out_valid),
    .io_data_1_out_bits(PE_199_io_data_1_out_bits),
    .io_data_0_in_valid(PE_199_io_data_0_in_valid),
    .io_data_0_in_bits(PE_199_io_data_0_in_bits),
    .io_data_0_out_valid(PE_199_io_data_0_out_valid),
    .io_data_0_out_bits(PE_199_io_data_0_out_bits)
  );
  PE PE_200 ( // @[pe.scala 187:13]
    .clock(PE_200_clock),
    .reset(PE_200_reset),
    .io_data_2_out_valid(PE_200_io_data_2_out_valid),
    .io_data_2_out_bits(PE_200_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_200_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_200_io_data_1_in_valid),
    .io_data_1_in_bits(PE_200_io_data_1_in_bits),
    .io_data_1_out_valid(PE_200_io_data_1_out_valid),
    .io_data_1_out_bits(PE_200_io_data_1_out_bits),
    .io_data_0_in_valid(PE_200_io_data_0_in_valid),
    .io_data_0_in_bits(PE_200_io_data_0_in_bits),
    .io_data_0_out_valid(PE_200_io_data_0_out_valid),
    .io_data_0_out_bits(PE_200_io_data_0_out_bits)
  );
  PE PE_201 ( // @[pe.scala 187:13]
    .clock(PE_201_clock),
    .reset(PE_201_reset),
    .io_data_2_out_valid(PE_201_io_data_2_out_valid),
    .io_data_2_out_bits(PE_201_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_201_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_201_io_data_1_in_valid),
    .io_data_1_in_bits(PE_201_io_data_1_in_bits),
    .io_data_1_out_valid(PE_201_io_data_1_out_valid),
    .io_data_1_out_bits(PE_201_io_data_1_out_bits),
    .io_data_0_in_valid(PE_201_io_data_0_in_valid),
    .io_data_0_in_bits(PE_201_io_data_0_in_bits),
    .io_data_0_out_valid(PE_201_io_data_0_out_valid),
    .io_data_0_out_bits(PE_201_io_data_0_out_bits)
  );
  PE PE_202 ( // @[pe.scala 187:13]
    .clock(PE_202_clock),
    .reset(PE_202_reset),
    .io_data_2_out_valid(PE_202_io_data_2_out_valid),
    .io_data_2_out_bits(PE_202_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_202_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_202_io_data_1_in_valid),
    .io_data_1_in_bits(PE_202_io_data_1_in_bits),
    .io_data_1_out_valid(PE_202_io_data_1_out_valid),
    .io_data_1_out_bits(PE_202_io_data_1_out_bits),
    .io_data_0_in_valid(PE_202_io_data_0_in_valid),
    .io_data_0_in_bits(PE_202_io_data_0_in_bits),
    .io_data_0_out_valid(PE_202_io_data_0_out_valid),
    .io_data_0_out_bits(PE_202_io_data_0_out_bits)
  );
  PE PE_203 ( // @[pe.scala 187:13]
    .clock(PE_203_clock),
    .reset(PE_203_reset),
    .io_data_2_out_valid(PE_203_io_data_2_out_valid),
    .io_data_2_out_bits(PE_203_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_203_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_203_io_data_1_in_valid),
    .io_data_1_in_bits(PE_203_io_data_1_in_bits),
    .io_data_1_out_valid(PE_203_io_data_1_out_valid),
    .io_data_1_out_bits(PE_203_io_data_1_out_bits),
    .io_data_0_in_valid(PE_203_io_data_0_in_valid),
    .io_data_0_in_bits(PE_203_io_data_0_in_bits),
    .io_data_0_out_valid(PE_203_io_data_0_out_valid),
    .io_data_0_out_bits(PE_203_io_data_0_out_bits)
  );
  PE PE_204 ( // @[pe.scala 187:13]
    .clock(PE_204_clock),
    .reset(PE_204_reset),
    .io_data_2_out_valid(PE_204_io_data_2_out_valid),
    .io_data_2_out_bits(PE_204_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_204_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_204_io_data_1_in_valid),
    .io_data_1_in_bits(PE_204_io_data_1_in_bits),
    .io_data_1_out_valid(PE_204_io_data_1_out_valid),
    .io_data_1_out_bits(PE_204_io_data_1_out_bits),
    .io_data_0_in_valid(PE_204_io_data_0_in_valid),
    .io_data_0_in_bits(PE_204_io_data_0_in_bits),
    .io_data_0_out_valid(PE_204_io_data_0_out_valid),
    .io_data_0_out_bits(PE_204_io_data_0_out_bits)
  );
  PE PE_205 ( // @[pe.scala 187:13]
    .clock(PE_205_clock),
    .reset(PE_205_reset),
    .io_data_2_out_valid(PE_205_io_data_2_out_valid),
    .io_data_2_out_bits(PE_205_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_205_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_205_io_data_1_in_valid),
    .io_data_1_in_bits(PE_205_io_data_1_in_bits),
    .io_data_1_out_valid(PE_205_io_data_1_out_valid),
    .io_data_1_out_bits(PE_205_io_data_1_out_bits),
    .io_data_0_in_valid(PE_205_io_data_0_in_valid),
    .io_data_0_in_bits(PE_205_io_data_0_in_bits),
    .io_data_0_out_valid(PE_205_io_data_0_out_valid),
    .io_data_0_out_bits(PE_205_io_data_0_out_bits)
  );
  PE PE_206 ( // @[pe.scala 187:13]
    .clock(PE_206_clock),
    .reset(PE_206_reset),
    .io_data_2_out_valid(PE_206_io_data_2_out_valid),
    .io_data_2_out_bits(PE_206_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_206_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_206_io_data_1_in_valid),
    .io_data_1_in_bits(PE_206_io_data_1_in_bits),
    .io_data_1_out_valid(PE_206_io_data_1_out_valid),
    .io_data_1_out_bits(PE_206_io_data_1_out_bits),
    .io_data_0_in_valid(PE_206_io_data_0_in_valid),
    .io_data_0_in_bits(PE_206_io_data_0_in_bits),
    .io_data_0_out_valid(PE_206_io_data_0_out_valid),
    .io_data_0_out_bits(PE_206_io_data_0_out_bits)
  );
  PE PE_207 ( // @[pe.scala 187:13]
    .clock(PE_207_clock),
    .reset(PE_207_reset),
    .io_data_2_out_valid(PE_207_io_data_2_out_valid),
    .io_data_2_out_bits(PE_207_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_207_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_207_io_data_1_in_valid),
    .io_data_1_in_bits(PE_207_io_data_1_in_bits),
    .io_data_1_out_valid(PE_207_io_data_1_out_valid),
    .io_data_1_out_bits(PE_207_io_data_1_out_bits),
    .io_data_0_in_valid(PE_207_io_data_0_in_valid),
    .io_data_0_in_bits(PE_207_io_data_0_in_bits),
    .io_data_0_out_valid(PE_207_io_data_0_out_valid),
    .io_data_0_out_bits(PE_207_io_data_0_out_bits)
  );
  PE PE_208 ( // @[pe.scala 187:13]
    .clock(PE_208_clock),
    .reset(PE_208_reset),
    .io_data_2_out_valid(PE_208_io_data_2_out_valid),
    .io_data_2_out_bits(PE_208_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_208_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_208_io_data_1_in_valid),
    .io_data_1_in_bits(PE_208_io_data_1_in_bits),
    .io_data_1_out_valid(PE_208_io_data_1_out_valid),
    .io_data_1_out_bits(PE_208_io_data_1_out_bits),
    .io_data_0_in_valid(PE_208_io_data_0_in_valid),
    .io_data_0_in_bits(PE_208_io_data_0_in_bits),
    .io_data_0_out_valid(PE_208_io_data_0_out_valid),
    .io_data_0_out_bits(PE_208_io_data_0_out_bits)
  );
  PE PE_209 ( // @[pe.scala 187:13]
    .clock(PE_209_clock),
    .reset(PE_209_reset),
    .io_data_2_out_valid(PE_209_io_data_2_out_valid),
    .io_data_2_out_bits(PE_209_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_209_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_209_io_data_1_in_valid),
    .io_data_1_in_bits(PE_209_io_data_1_in_bits),
    .io_data_1_out_valid(PE_209_io_data_1_out_valid),
    .io_data_1_out_bits(PE_209_io_data_1_out_bits),
    .io_data_0_in_valid(PE_209_io_data_0_in_valid),
    .io_data_0_in_bits(PE_209_io_data_0_in_bits),
    .io_data_0_out_valid(PE_209_io_data_0_out_valid),
    .io_data_0_out_bits(PE_209_io_data_0_out_bits)
  );
  PE PE_210 ( // @[pe.scala 187:13]
    .clock(PE_210_clock),
    .reset(PE_210_reset),
    .io_data_2_out_valid(PE_210_io_data_2_out_valid),
    .io_data_2_out_bits(PE_210_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_210_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_210_io_data_1_in_valid),
    .io_data_1_in_bits(PE_210_io_data_1_in_bits),
    .io_data_1_out_valid(PE_210_io_data_1_out_valid),
    .io_data_1_out_bits(PE_210_io_data_1_out_bits),
    .io_data_0_in_valid(PE_210_io_data_0_in_valid),
    .io_data_0_in_bits(PE_210_io_data_0_in_bits),
    .io_data_0_out_valid(PE_210_io_data_0_out_valid),
    .io_data_0_out_bits(PE_210_io_data_0_out_bits)
  );
  PE PE_211 ( // @[pe.scala 187:13]
    .clock(PE_211_clock),
    .reset(PE_211_reset),
    .io_data_2_out_valid(PE_211_io_data_2_out_valid),
    .io_data_2_out_bits(PE_211_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_211_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_211_io_data_1_in_valid),
    .io_data_1_in_bits(PE_211_io_data_1_in_bits),
    .io_data_1_out_valid(PE_211_io_data_1_out_valid),
    .io_data_1_out_bits(PE_211_io_data_1_out_bits),
    .io_data_0_in_valid(PE_211_io_data_0_in_valid),
    .io_data_0_in_bits(PE_211_io_data_0_in_bits),
    .io_data_0_out_valid(PE_211_io_data_0_out_valid),
    .io_data_0_out_bits(PE_211_io_data_0_out_bits)
  );
  PE PE_212 ( // @[pe.scala 187:13]
    .clock(PE_212_clock),
    .reset(PE_212_reset),
    .io_data_2_out_valid(PE_212_io_data_2_out_valid),
    .io_data_2_out_bits(PE_212_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_212_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_212_io_data_1_in_valid),
    .io_data_1_in_bits(PE_212_io_data_1_in_bits),
    .io_data_1_out_valid(PE_212_io_data_1_out_valid),
    .io_data_1_out_bits(PE_212_io_data_1_out_bits),
    .io_data_0_in_valid(PE_212_io_data_0_in_valid),
    .io_data_0_in_bits(PE_212_io_data_0_in_bits),
    .io_data_0_out_valid(PE_212_io_data_0_out_valid),
    .io_data_0_out_bits(PE_212_io_data_0_out_bits)
  );
  PE PE_213 ( // @[pe.scala 187:13]
    .clock(PE_213_clock),
    .reset(PE_213_reset),
    .io_data_2_out_valid(PE_213_io_data_2_out_valid),
    .io_data_2_out_bits(PE_213_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_213_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_213_io_data_1_in_valid),
    .io_data_1_in_bits(PE_213_io_data_1_in_bits),
    .io_data_1_out_valid(PE_213_io_data_1_out_valid),
    .io_data_1_out_bits(PE_213_io_data_1_out_bits),
    .io_data_0_in_valid(PE_213_io_data_0_in_valid),
    .io_data_0_in_bits(PE_213_io_data_0_in_bits),
    .io_data_0_out_valid(PE_213_io_data_0_out_valid),
    .io_data_0_out_bits(PE_213_io_data_0_out_bits)
  );
  PE PE_214 ( // @[pe.scala 187:13]
    .clock(PE_214_clock),
    .reset(PE_214_reset),
    .io_data_2_out_valid(PE_214_io_data_2_out_valid),
    .io_data_2_out_bits(PE_214_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_214_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_214_io_data_1_in_valid),
    .io_data_1_in_bits(PE_214_io_data_1_in_bits),
    .io_data_1_out_valid(PE_214_io_data_1_out_valid),
    .io_data_1_out_bits(PE_214_io_data_1_out_bits),
    .io_data_0_in_valid(PE_214_io_data_0_in_valid),
    .io_data_0_in_bits(PE_214_io_data_0_in_bits),
    .io_data_0_out_valid(PE_214_io_data_0_out_valid),
    .io_data_0_out_bits(PE_214_io_data_0_out_bits)
  );
  PE PE_215 ( // @[pe.scala 187:13]
    .clock(PE_215_clock),
    .reset(PE_215_reset),
    .io_data_2_out_valid(PE_215_io_data_2_out_valid),
    .io_data_2_out_bits(PE_215_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_215_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_215_io_data_1_in_valid),
    .io_data_1_in_bits(PE_215_io_data_1_in_bits),
    .io_data_1_out_valid(PE_215_io_data_1_out_valid),
    .io_data_1_out_bits(PE_215_io_data_1_out_bits),
    .io_data_0_in_valid(PE_215_io_data_0_in_valid),
    .io_data_0_in_bits(PE_215_io_data_0_in_bits),
    .io_data_0_out_valid(PE_215_io_data_0_out_valid),
    .io_data_0_out_bits(PE_215_io_data_0_out_bits)
  );
  PE PE_216 ( // @[pe.scala 187:13]
    .clock(PE_216_clock),
    .reset(PE_216_reset),
    .io_data_2_out_valid(PE_216_io_data_2_out_valid),
    .io_data_2_out_bits(PE_216_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_216_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_216_io_data_1_in_valid),
    .io_data_1_in_bits(PE_216_io_data_1_in_bits),
    .io_data_1_out_valid(PE_216_io_data_1_out_valid),
    .io_data_1_out_bits(PE_216_io_data_1_out_bits),
    .io_data_0_in_valid(PE_216_io_data_0_in_valid),
    .io_data_0_in_bits(PE_216_io_data_0_in_bits),
    .io_data_0_out_valid(PE_216_io_data_0_out_valid),
    .io_data_0_out_bits(PE_216_io_data_0_out_bits)
  );
  PE PE_217 ( // @[pe.scala 187:13]
    .clock(PE_217_clock),
    .reset(PE_217_reset),
    .io_data_2_out_valid(PE_217_io_data_2_out_valid),
    .io_data_2_out_bits(PE_217_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_217_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_217_io_data_1_in_valid),
    .io_data_1_in_bits(PE_217_io_data_1_in_bits),
    .io_data_1_out_valid(PE_217_io_data_1_out_valid),
    .io_data_1_out_bits(PE_217_io_data_1_out_bits),
    .io_data_0_in_valid(PE_217_io_data_0_in_valid),
    .io_data_0_in_bits(PE_217_io_data_0_in_bits),
    .io_data_0_out_valid(PE_217_io_data_0_out_valid),
    .io_data_0_out_bits(PE_217_io_data_0_out_bits)
  );
  PE PE_218 ( // @[pe.scala 187:13]
    .clock(PE_218_clock),
    .reset(PE_218_reset),
    .io_data_2_out_valid(PE_218_io_data_2_out_valid),
    .io_data_2_out_bits(PE_218_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_218_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_218_io_data_1_in_valid),
    .io_data_1_in_bits(PE_218_io_data_1_in_bits),
    .io_data_1_out_valid(PE_218_io_data_1_out_valid),
    .io_data_1_out_bits(PE_218_io_data_1_out_bits),
    .io_data_0_in_valid(PE_218_io_data_0_in_valid),
    .io_data_0_in_bits(PE_218_io_data_0_in_bits),
    .io_data_0_out_valid(PE_218_io_data_0_out_valid),
    .io_data_0_out_bits(PE_218_io_data_0_out_bits)
  );
  PE PE_219 ( // @[pe.scala 187:13]
    .clock(PE_219_clock),
    .reset(PE_219_reset),
    .io_data_2_out_valid(PE_219_io_data_2_out_valid),
    .io_data_2_out_bits(PE_219_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_219_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_219_io_data_1_in_valid),
    .io_data_1_in_bits(PE_219_io_data_1_in_bits),
    .io_data_1_out_valid(PE_219_io_data_1_out_valid),
    .io_data_1_out_bits(PE_219_io_data_1_out_bits),
    .io_data_0_in_valid(PE_219_io_data_0_in_valid),
    .io_data_0_in_bits(PE_219_io_data_0_in_bits),
    .io_data_0_out_valid(PE_219_io_data_0_out_valid),
    .io_data_0_out_bits(PE_219_io_data_0_out_bits)
  );
  PE PE_220 ( // @[pe.scala 187:13]
    .clock(PE_220_clock),
    .reset(PE_220_reset),
    .io_data_2_out_valid(PE_220_io_data_2_out_valid),
    .io_data_2_out_bits(PE_220_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_220_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_220_io_data_1_in_valid),
    .io_data_1_in_bits(PE_220_io_data_1_in_bits),
    .io_data_1_out_valid(PE_220_io_data_1_out_valid),
    .io_data_1_out_bits(PE_220_io_data_1_out_bits),
    .io_data_0_in_valid(PE_220_io_data_0_in_valid),
    .io_data_0_in_bits(PE_220_io_data_0_in_bits),
    .io_data_0_out_valid(PE_220_io_data_0_out_valid),
    .io_data_0_out_bits(PE_220_io_data_0_out_bits)
  );
  PE PE_221 ( // @[pe.scala 187:13]
    .clock(PE_221_clock),
    .reset(PE_221_reset),
    .io_data_2_out_valid(PE_221_io_data_2_out_valid),
    .io_data_2_out_bits(PE_221_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_221_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_221_io_data_1_in_valid),
    .io_data_1_in_bits(PE_221_io_data_1_in_bits),
    .io_data_1_out_valid(PE_221_io_data_1_out_valid),
    .io_data_1_out_bits(PE_221_io_data_1_out_bits),
    .io_data_0_in_valid(PE_221_io_data_0_in_valid),
    .io_data_0_in_bits(PE_221_io_data_0_in_bits),
    .io_data_0_out_valid(PE_221_io_data_0_out_valid),
    .io_data_0_out_bits(PE_221_io_data_0_out_bits)
  );
  PE PE_222 ( // @[pe.scala 187:13]
    .clock(PE_222_clock),
    .reset(PE_222_reset),
    .io_data_2_out_valid(PE_222_io_data_2_out_valid),
    .io_data_2_out_bits(PE_222_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_222_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_222_io_data_1_in_valid),
    .io_data_1_in_bits(PE_222_io_data_1_in_bits),
    .io_data_1_out_valid(PE_222_io_data_1_out_valid),
    .io_data_1_out_bits(PE_222_io_data_1_out_bits),
    .io_data_0_in_valid(PE_222_io_data_0_in_valid),
    .io_data_0_in_bits(PE_222_io_data_0_in_bits),
    .io_data_0_out_valid(PE_222_io_data_0_out_valid),
    .io_data_0_out_bits(PE_222_io_data_0_out_bits)
  );
  PE PE_223 ( // @[pe.scala 187:13]
    .clock(PE_223_clock),
    .reset(PE_223_reset),
    .io_data_2_out_valid(PE_223_io_data_2_out_valid),
    .io_data_2_out_bits(PE_223_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_223_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_223_io_data_1_in_valid),
    .io_data_1_in_bits(PE_223_io_data_1_in_bits),
    .io_data_1_out_valid(PE_223_io_data_1_out_valid),
    .io_data_1_out_bits(PE_223_io_data_1_out_bits),
    .io_data_0_in_valid(PE_223_io_data_0_in_valid),
    .io_data_0_in_bits(PE_223_io_data_0_in_bits),
    .io_data_0_out_valid(PE_223_io_data_0_out_valid),
    .io_data_0_out_bits(PE_223_io_data_0_out_bits)
  );
  PE PE_224 ( // @[pe.scala 187:13]
    .clock(PE_224_clock),
    .reset(PE_224_reset),
    .io_data_2_out_valid(PE_224_io_data_2_out_valid),
    .io_data_2_out_bits(PE_224_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_224_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_224_io_data_1_in_valid),
    .io_data_1_in_bits(PE_224_io_data_1_in_bits),
    .io_data_1_out_valid(PE_224_io_data_1_out_valid),
    .io_data_1_out_bits(PE_224_io_data_1_out_bits),
    .io_data_0_in_valid(PE_224_io_data_0_in_valid),
    .io_data_0_in_bits(PE_224_io_data_0_in_bits),
    .io_data_0_out_valid(PE_224_io_data_0_out_valid),
    .io_data_0_out_bits(PE_224_io_data_0_out_bits)
  );
  PE PE_225 ( // @[pe.scala 187:13]
    .clock(PE_225_clock),
    .reset(PE_225_reset),
    .io_data_2_out_valid(PE_225_io_data_2_out_valid),
    .io_data_2_out_bits(PE_225_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_225_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_225_io_data_1_in_valid),
    .io_data_1_in_bits(PE_225_io_data_1_in_bits),
    .io_data_1_out_valid(PE_225_io_data_1_out_valid),
    .io_data_1_out_bits(PE_225_io_data_1_out_bits),
    .io_data_0_in_valid(PE_225_io_data_0_in_valid),
    .io_data_0_in_bits(PE_225_io_data_0_in_bits),
    .io_data_0_out_valid(PE_225_io_data_0_out_valid),
    .io_data_0_out_bits(PE_225_io_data_0_out_bits)
  );
  PE PE_226 ( // @[pe.scala 187:13]
    .clock(PE_226_clock),
    .reset(PE_226_reset),
    .io_data_2_out_valid(PE_226_io_data_2_out_valid),
    .io_data_2_out_bits(PE_226_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_226_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_226_io_data_1_in_valid),
    .io_data_1_in_bits(PE_226_io_data_1_in_bits),
    .io_data_1_out_valid(PE_226_io_data_1_out_valid),
    .io_data_1_out_bits(PE_226_io_data_1_out_bits),
    .io_data_0_in_valid(PE_226_io_data_0_in_valid),
    .io_data_0_in_bits(PE_226_io_data_0_in_bits),
    .io_data_0_out_valid(PE_226_io_data_0_out_valid),
    .io_data_0_out_bits(PE_226_io_data_0_out_bits)
  );
  PE PE_227 ( // @[pe.scala 187:13]
    .clock(PE_227_clock),
    .reset(PE_227_reset),
    .io_data_2_out_valid(PE_227_io_data_2_out_valid),
    .io_data_2_out_bits(PE_227_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_227_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_227_io_data_1_in_valid),
    .io_data_1_in_bits(PE_227_io_data_1_in_bits),
    .io_data_1_out_valid(PE_227_io_data_1_out_valid),
    .io_data_1_out_bits(PE_227_io_data_1_out_bits),
    .io_data_0_in_valid(PE_227_io_data_0_in_valid),
    .io_data_0_in_bits(PE_227_io_data_0_in_bits),
    .io_data_0_out_valid(PE_227_io_data_0_out_valid),
    .io_data_0_out_bits(PE_227_io_data_0_out_bits)
  );
  PE PE_228 ( // @[pe.scala 187:13]
    .clock(PE_228_clock),
    .reset(PE_228_reset),
    .io_data_2_out_valid(PE_228_io_data_2_out_valid),
    .io_data_2_out_bits(PE_228_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_228_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_228_io_data_1_in_valid),
    .io_data_1_in_bits(PE_228_io_data_1_in_bits),
    .io_data_1_out_valid(PE_228_io_data_1_out_valid),
    .io_data_1_out_bits(PE_228_io_data_1_out_bits),
    .io_data_0_in_valid(PE_228_io_data_0_in_valid),
    .io_data_0_in_bits(PE_228_io_data_0_in_bits),
    .io_data_0_out_valid(PE_228_io_data_0_out_valid),
    .io_data_0_out_bits(PE_228_io_data_0_out_bits)
  );
  PE PE_229 ( // @[pe.scala 187:13]
    .clock(PE_229_clock),
    .reset(PE_229_reset),
    .io_data_2_out_valid(PE_229_io_data_2_out_valid),
    .io_data_2_out_bits(PE_229_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_229_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_229_io_data_1_in_valid),
    .io_data_1_in_bits(PE_229_io_data_1_in_bits),
    .io_data_1_out_valid(PE_229_io_data_1_out_valid),
    .io_data_1_out_bits(PE_229_io_data_1_out_bits),
    .io_data_0_in_valid(PE_229_io_data_0_in_valid),
    .io_data_0_in_bits(PE_229_io_data_0_in_bits),
    .io_data_0_out_valid(PE_229_io_data_0_out_valid),
    .io_data_0_out_bits(PE_229_io_data_0_out_bits)
  );
  PE PE_230 ( // @[pe.scala 187:13]
    .clock(PE_230_clock),
    .reset(PE_230_reset),
    .io_data_2_out_valid(PE_230_io_data_2_out_valid),
    .io_data_2_out_bits(PE_230_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_230_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_230_io_data_1_in_valid),
    .io_data_1_in_bits(PE_230_io_data_1_in_bits),
    .io_data_1_out_valid(PE_230_io_data_1_out_valid),
    .io_data_1_out_bits(PE_230_io_data_1_out_bits),
    .io_data_0_in_valid(PE_230_io_data_0_in_valid),
    .io_data_0_in_bits(PE_230_io_data_0_in_bits),
    .io_data_0_out_valid(PE_230_io_data_0_out_valid),
    .io_data_0_out_bits(PE_230_io_data_0_out_bits)
  );
  PE PE_231 ( // @[pe.scala 187:13]
    .clock(PE_231_clock),
    .reset(PE_231_reset),
    .io_data_2_out_valid(PE_231_io_data_2_out_valid),
    .io_data_2_out_bits(PE_231_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_231_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_231_io_data_1_in_valid),
    .io_data_1_in_bits(PE_231_io_data_1_in_bits),
    .io_data_1_out_valid(PE_231_io_data_1_out_valid),
    .io_data_1_out_bits(PE_231_io_data_1_out_bits),
    .io_data_0_in_valid(PE_231_io_data_0_in_valid),
    .io_data_0_in_bits(PE_231_io_data_0_in_bits),
    .io_data_0_out_valid(PE_231_io_data_0_out_valid),
    .io_data_0_out_bits(PE_231_io_data_0_out_bits)
  );
  PE PE_232 ( // @[pe.scala 187:13]
    .clock(PE_232_clock),
    .reset(PE_232_reset),
    .io_data_2_out_valid(PE_232_io_data_2_out_valid),
    .io_data_2_out_bits(PE_232_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_232_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_232_io_data_1_in_valid),
    .io_data_1_in_bits(PE_232_io_data_1_in_bits),
    .io_data_1_out_valid(PE_232_io_data_1_out_valid),
    .io_data_1_out_bits(PE_232_io_data_1_out_bits),
    .io_data_0_in_valid(PE_232_io_data_0_in_valid),
    .io_data_0_in_bits(PE_232_io_data_0_in_bits),
    .io_data_0_out_valid(PE_232_io_data_0_out_valid),
    .io_data_0_out_bits(PE_232_io_data_0_out_bits)
  );
  PE PE_233 ( // @[pe.scala 187:13]
    .clock(PE_233_clock),
    .reset(PE_233_reset),
    .io_data_2_out_valid(PE_233_io_data_2_out_valid),
    .io_data_2_out_bits(PE_233_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_233_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_233_io_data_1_in_valid),
    .io_data_1_in_bits(PE_233_io_data_1_in_bits),
    .io_data_1_out_valid(PE_233_io_data_1_out_valid),
    .io_data_1_out_bits(PE_233_io_data_1_out_bits),
    .io_data_0_in_valid(PE_233_io_data_0_in_valid),
    .io_data_0_in_bits(PE_233_io_data_0_in_bits),
    .io_data_0_out_valid(PE_233_io_data_0_out_valid),
    .io_data_0_out_bits(PE_233_io_data_0_out_bits)
  );
  PE PE_234 ( // @[pe.scala 187:13]
    .clock(PE_234_clock),
    .reset(PE_234_reset),
    .io_data_2_out_valid(PE_234_io_data_2_out_valid),
    .io_data_2_out_bits(PE_234_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_234_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_234_io_data_1_in_valid),
    .io_data_1_in_bits(PE_234_io_data_1_in_bits),
    .io_data_1_out_valid(PE_234_io_data_1_out_valid),
    .io_data_1_out_bits(PE_234_io_data_1_out_bits),
    .io_data_0_in_valid(PE_234_io_data_0_in_valid),
    .io_data_0_in_bits(PE_234_io_data_0_in_bits),
    .io_data_0_out_valid(PE_234_io_data_0_out_valid),
    .io_data_0_out_bits(PE_234_io_data_0_out_bits)
  );
  PE PE_235 ( // @[pe.scala 187:13]
    .clock(PE_235_clock),
    .reset(PE_235_reset),
    .io_data_2_out_valid(PE_235_io_data_2_out_valid),
    .io_data_2_out_bits(PE_235_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_235_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_235_io_data_1_in_valid),
    .io_data_1_in_bits(PE_235_io_data_1_in_bits),
    .io_data_1_out_valid(PE_235_io_data_1_out_valid),
    .io_data_1_out_bits(PE_235_io_data_1_out_bits),
    .io_data_0_in_valid(PE_235_io_data_0_in_valid),
    .io_data_0_in_bits(PE_235_io_data_0_in_bits),
    .io_data_0_out_valid(PE_235_io_data_0_out_valid),
    .io_data_0_out_bits(PE_235_io_data_0_out_bits)
  );
  PE PE_236 ( // @[pe.scala 187:13]
    .clock(PE_236_clock),
    .reset(PE_236_reset),
    .io_data_2_out_valid(PE_236_io_data_2_out_valid),
    .io_data_2_out_bits(PE_236_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_236_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_236_io_data_1_in_valid),
    .io_data_1_in_bits(PE_236_io_data_1_in_bits),
    .io_data_1_out_valid(PE_236_io_data_1_out_valid),
    .io_data_1_out_bits(PE_236_io_data_1_out_bits),
    .io_data_0_in_valid(PE_236_io_data_0_in_valid),
    .io_data_0_in_bits(PE_236_io_data_0_in_bits),
    .io_data_0_out_valid(PE_236_io_data_0_out_valid),
    .io_data_0_out_bits(PE_236_io_data_0_out_bits)
  );
  PE PE_237 ( // @[pe.scala 187:13]
    .clock(PE_237_clock),
    .reset(PE_237_reset),
    .io_data_2_out_valid(PE_237_io_data_2_out_valid),
    .io_data_2_out_bits(PE_237_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_237_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_237_io_data_1_in_valid),
    .io_data_1_in_bits(PE_237_io_data_1_in_bits),
    .io_data_1_out_valid(PE_237_io_data_1_out_valid),
    .io_data_1_out_bits(PE_237_io_data_1_out_bits),
    .io_data_0_in_valid(PE_237_io_data_0_in_valid),
    .io_data_0_in_bits(PE_237_io_data_0_in_bits),
    .io_data_0_out_valid(PE_237_io_data_0_out_valid),
    .io_data_0_out_bits(PE_237_io_data_0_out_bits)
  );
  PE PE_238 ( // @[pe.scala 187:13]
    .clock(PE_238_clock),
    .reset(PE_238_reset),
    .io_data_2_out_valid(PE_238_io_data_2_out_valid),
    .io_data_2_out_bits(PE_238_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_238_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_238_io_data_1_in_valid),
    .io_data_1_in_bits(PE_238_io_data_1_in_bits),
    .io_data_1_out_valid(PE_238_io_data_1_out_valid),
    .io_data_1_out_bits(PE_238_io_data_1_out_bits),
    .io_data_0_in_valid(PE_238_io_data_0_in_valid),
    .io_data_0_in_bits(PE_238_io_data_0_in_bits),
    .io_data_0_out_valid(PE_238_io_data_0_out_valid),
    .io_data_0_out_bits(PE_238_io_data_0_out_bits)
  );
  PE PE_239 ( // @[pe.scala 187:13]
    .clock(PE_239_clock),
    .reset(PE_239_reset),
    .io_data_2_out_valid(PE_239_io_data_2_out_valid),
    .io_data_2_out_bits(PE_239_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_239_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_239_io_data_1_in_valid),
    .io_data_1_in_bits(PE_239_io_data_1_in_bits),
    .io_data_1_out_valid(PE_239_io_data_1_out_valid),
    .io_data_1_out_bits(PE_239_io_data_1_out_bits),
    .io_data_0_in_valid(PE_239_io_data_0_in_valid),
    .io_data_0_in_bits(PE_239_io_data_0_in_bits),
    .io_data_0_out_valid(PE_239_io_data_0_out_valid),
    .io_data_0_out_bits(PE_239_io_data_0_out_bits)
  );
  PE PE_240 ( // @[pe.scala 187:13]
    .clock(PE_240_clock),
    .reset(PE_240_reset),
    .io_data_2_out_valid(PE_240_io_data_2_out_valid),
    .io_data_2_out_bits(PE_240_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_240_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_240_io_data_1_in_valid),
    .io_data_1_in_bits(PE_240_io_data_1_in_bits),
    .io_data_1_out_valid(PE_240_io_data_1_out_valid),
    .io_data_1_out_bits(PE_240_io_data_1_out_bits),
    .io_data_0_in_valid(PE_240_io_data_0_in_valid),
    .io_data_0_in_bits(PE_240_io_data_0_in_bits),
    .io_data_0_out_valid(PE_240_io_data_0_out_valid),
    .io_data_0_out_bits(PE_240_io_data_0_out_bits)
  );
  PE PE_241 ( // @[pe.scala 187:13]
    .clock(PE_241_clock),
    .reset(PE_241_reset),
    .io_data_2_out_valid(PE_241_io_data_2_out_valid),
    .io_data_2_out_bits(PE_241_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_241_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_241_io_data_1_in_valid),
    .io_data_1_in_bits(PE_241_io_data_1_in_bits),
    .io_data_1_out_valid(PE_241_io_data_1_out_valid),
    .io_data_1_out_bits(PE_241_io_data_1_out_bits),
    .io_data_0_in_valid(PE_241_io_data_0_in_valid),
    .io_data_0_in_bits(PE_241_io_data_0_in_bits),
    .io_data_0_out_valid(PE_241_io_data_0_out_valid),
    .io_data_0_out_bits(PE_241_io_data_0_out_bits)
  );
  PE PE_242 ( // @[pe.scala 187:13]
    .clock(PE_242_clock),
    .reset(PE_242_reset),
    .io_data_2_out_valid(PE_242_io_data_2_out_valid),
    .io_data_2_out_bits(PE_242_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_242_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_242_io_data_1_in_valid),
    .io_data_1_in_bits(PE_242_io_data_1_in_bits),
    .io_data_1_out_valid(PE_242_io_data_1_out_valid),
    .io_data_1_out_bits(PE_242_io_data_1_out_bits),
    .io_data_0_in_valid(PE_242_io_data_0_in_valid),
    .io_data_0_in_bits(PE_242_io_data_0_in_bits),
    .io_data_0_out_valid(PE_242_io_data_0_out_valid),
    .io_data_0_out_bits(PE_242_io_data_0_out_bits)
  );
  PE PE_243 ( // @[pe.scala 187:13]
    .clock(PE_243_clock),
    .reset(PE_243_reset),
    .io_data_2_out_valid(PE_243_io_data_2_out_valid),
    .io_data_2_out_bits(PE_243_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_243_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_243_io_data_1_in_valid),
    .io_data_1_in_bits(PE_243_io_data_1_in_bits),
    .io_data_1_out_valid(PE_243_io_data_1_out_valid),
    .io_data_1_out_bits(PE_243_io_data_1_out_bits),
    .io_data_0_in_valid(PE_243_io_data_0_in_valid),
    .io_data_0_in_bits(PE_243_io_data_0_in_bits),
    .io_data_0_out_valid(PE_243_io_data_0_out_valid),
    .io_data_0_out_bits(PE_243_io_data_0_out_bits)
  );
  PE PE_244 ( // @[pe.scala 187:13]
    .clock(PE_244_clock),
    .reset(PE_244_reset),
    .io_data_2_out_valid(PE_244_io_data_2_out_valid),
    .io_data_2_out_bits(PE_244_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_244_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_244_io_data_1_in_valid),
    .io_data_1_in_bits(PE_244_io_data_1_in_bits),
    .io_data_1_out_valid(PE_244_io_data_1_out_valid),
    .io_data_1_out_bits(PE_244_io_data_1_out_bits),
    .io_data_0_in_valid(PE_244_io_data_0_in_valid),
    .io_data_0_in_bits(PE_244_io_data_0_in_bits),
    .io_data_0_out_valid(PE_244_io_data_0_out_valid),
    .io_data_0_out_bits(PE_244_io_data_0_out_bits)
  );
  PE PE_245 ( // @[pe.scala 187:13]
    .clock(PE_245_clock),
    .reset(PE_245_reset),
    .io_data_2_out_valid(PE_245_io_data_2_out_valid),
    .io_data_2_out_bits(PE_245_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_245_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_245_io_data_1_in_valid),
    .io_data_1_in_bits(PE_245_io_data_1_in_bits),
    .io_data_1_out_valid(PE_245_io_data_1_out_valid),
    .io_data_1_out_bits(PE_245_io_data_1_out_bits),
    .io_data_0_in_valid(PE_245_io_data_0_in_valid),
    .io_data_0_in_bits(PE_245_io_data_0_in_bits),
    .io_data_0_out_valid(PE_245_io_data_0_out_valid),
    .io_data_0_out_bits(PE_245_io_data_0_out_bits)
  );
  PE PE_246 ( // @[pe.scala 187:13]
    .clock(PE_246_clock),
    .reset(PE_246_reset),
    .io_data_2_out_valid(PE_246_io_data_2_out_valid),
    .io_data_2_out_bits(PE_246_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_246_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_246_io_data_1_in_valid),
    .io_data_1_in_bits(PE_246_io_data_1_in_bits),
    .io_data_1_out_valid(PE_246_io_data_1_out_valid),
    .io_data_1_out_bits(PE_246_io_data_1_out_bits),
    .io_data_0_in_valid(PE_246_io_data_0_in_valid),
    .io_data_0_in_bits(PE_246_io_data_0_in_bits),
    .io_data_0_out_valid(PE_246_io_data_0_out_valid),
    .io_data_0_out_bits(PE_246_io_data_0_out_bits)
  );
  PE PE_247 ( // @[pe.scala 187:13]
    .clock(PE_247_clock),
    .reset(PE_247_reset),
    .io_data_2_out_valid(PE_247_io_data_2_out_valid),
    .io_data_2_out_bits(PE_247_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_247_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_247_io_data_1_in_valid),
    .io_data_1_in_bits(PE_247_io_data_1_in_bits),
    .io_data_1_out_valid(PE_247_io_data_1_out_valid),
    .io_data_1_out_bits(PE_247_io_data_1_out_bits),
    .io_data_0_in_valid(PE_247_io_data_0_in_valid),
    .io_data_0_in_bits(PE_247_io_data_0_in_bits),
    .io_data_0_out_valid(PE_247_io_data_0_out_valid),
    .io_data_0_out_bits(PE_247_io_data_0_out_bits)
  );
  PE PE_248 ( // @[pe.scala 187:13]
    .clock(PE_248_clock),
    .reset(PE_248_reset),
    .io_data_2_out_valid(PE_248_io_data_2_out_valid),
    .io_data_2_out_bits(PE_248_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_248_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_248_io_data_1_in_valid),
    .io_data_1_in_bits(PE_248_io_data_1_in_bits),
    .io_data_1_out_valid(PE_248_io_data_1_out_valid),
    .io_data_1_out_bits(PE_248_io_data_1_out_bits),
    .io_data_0_in_valid(PE_248_io_data_0_in_valid),
    .io_data_0_in_bits(PE_248_io_data_0_in_bits),
    .io_data_0_out_valid(PE_248_io_data_0_out_valid),
    .io_data_0_out_bits(PE_248_io_data_0_out_bits)
  );
  PE PE_249 ( // @[pe.scala 187:13]
    .clock(PE_249_clock),
    .reset(PE_249_reset),
    .io_data_2_out_valid(PE_249_io_data_2_out_valid),
    .io_data_2_out_bits(PE_249_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_249_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_249_io_data_1_in_valid),
    .io_data_1_in_bits(PE_249_io_data_1_in_bits),
    .io_data_1_out_valid(PE_249_io_data_1_out_valid),
    .io_data_1_out_bits(PE_249_io_data_1_out_bits),
    .io_data_0_in_valid(PE_249_io_data_0_in_valid),
    .io_data_0_in_bits(PE_249_io_data_0_in_bits),
    .io_data_0_out_valid(PE_249_io_data_0_out_valid),
    .io_data_0_out_bits(PE_249_io_data_0_out_bits)
  );
  PE PE_250 ( // @[pe.scala 187:13]
    .clock(PE_250_clock),
    .reset(PE_250_reset),
    .io_data_2_out_valid(PE_250_io_data_2_out_valid),
    .io_data_2_out_bits(PE_250_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_250_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_250_io_data_1_in_valid),
    .io_data_1_in_bits(PE_250_io_data_1_in_bits),
    .io_data_1_out_valid(PE_250_io_data_1_out_valid),
    .io_data_1_out_bits(PE_250_io_data_1_out_bits),
    .io_data_0_in_valid(PE_250_io_data_0_in_valid),
    .io_data_0_in_bits(PE_250_io_data_0_in_bits),
    .io_data_0_out_valid(PE_250_io_data_0_out_valid),
    .io_data_0_out_bits(PE_250_io_data_0_out_bits)
  );
  PE PE_251 ( // @[pe.scala 187:13]
    .clock(PE_251_clock),
    .reset(PE_251_reset),
    .io_data_2_out_valid(PE_251_io_data_2_out_valid),
    .io_data_2_out_bits(PE_251_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_251_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_251_io_data_1_in_valid),
    .io_data_1_in_bits(PE_251_io_data_1_in_bits),
    .io_data_1_out_valid(PE_251_io_data_1_out_valid),
    .io_data_1_out_bits(PE_251_io_data_1_out_bits),
    .io_data_0_in_valid(PE_251_io_data_0_in_valid),
    .io_data_0_in_bits(PE_251_io_data_0_in_bits),
    .io_data_0_out_valid(PE_251_io_data_0_out_valid),
    .io_data_0_out_bits(PE_251_io_data_0_out_bits)
  );
  PE PE_252 ( // @[pe.scala 187:13]
    .clock(PE_252_clock),
    .reset(PE_252_reset),
    .io_data_2_out_valid(PE_252_io_data_2_out_valid),
    .io_data_2_out_bits(PE_252_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_252_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_252_io_data_1_in_valid),
    .io_data_1_in_bits(PE_252_io_data_1_in_bits),
    .io_data_1_out_valid(PE_252_io_data_1_out_valid),
    .io_data_1_out_bits(PE_252_io_data_1_out_bits),
    .io_data_0_in_valid(PE_252_io_data_0_in_valid),
    .io_data_0_in_bits(PE_252_io_data_0_in_bits),
    .io_data_0_out_valid(PE_252_io_data_0_out_valid),
    .io_data_0_out_bits(PE_252_io_data_0_out_bits)
  );
  PE PE_253 ( // @[pe.scala 187:13]
    .clock(PE_253_clock),
    .reset(PE_253_reset),
    .io_data_2_out_valid(PE_253_io_data_2_out_valid),
    .io_data_2_out_bits(PE_253_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_253_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_253_io_data_1_in_valid),
    .io_data_1_in_bits(PE_253_io_data_1_in_bits),
    .io_data_1_out_valid(PE_253_io_data_1_out_valid),
    .io_data_1_out_bits(PE_253_io_data_1_out_bits),
    .io_data_0_in_valid(PE_253_io_data_0_in_valid),
    .io_data_0_in_bits(PE_253_io_data_0_in_bits),
    .io_data_0_out_valid(PE_253_io_data_0_out_valid),
    .io_data_0_out_bits(PE_253_io_data_0_out_bits)
  );
  PE PE_254 ( // @[pe.scala 187:13]
    .clock(PE_254_clock),
    .reset(PE_254_reset),
    .io_data_2_out_valid(PE_254_io_data_2_out_valid),
    .io_data_2_out_bits(PE_254_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_254_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_254_io_data_1_in_valid),
    .io_data_1_in_bits(PE_254_io_data_1_in_bits),
    .io_data_1_out_valid(PE_254_io_data_1_out_valid),
    .io_data_1_out_bits(PE_254_io_data_1_out_bits),
    .io_data_0_in_valid(PE_254_io_data_0_in_valid),
    .io_data_0_in_bits(PE_254_io_data_0_in_bits),
    .io_data_0_out_valid(PE_254_io_data_0_out_valid),
    .io_data_0_out_bits(PE_254_io_data_0_out_bits)
  );
  PE PE_255 ( // @[pe.scala 187:13]
    .clock(PE_255_clock),
    .reset(PE_255_reset),
    .io_data_2_out_valid(PE_255_io_data_2_out_valid),
    .io_data_2_out_bits(PE_255_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_255_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_255_io_data_1_in_valid),
    .io_data_1_in_bits(PE_255_io_data_1_in_bits),
    .io_data_1_out_valid(PE_255_io_data_1_out_valid),
    .io_data_1_out_bits(PE_255_io_data_1_out_bits),
    .io_data_0_in_valid(PE_255_io_data_0_in_valid),
    .io_data_0_in_bits(PE_255_io_data_0_in_bits),
    .io_data_0_out_valid(PE_255_io_data_0_out_valid),
    .io_data_0_out_bits(PE_255_io_data_0_out_bits)
  );
  PE PE_256 ( // @[pe.scala 187:13]
    .clock(PE_256_clock),
    .reset(PE_256_reset),
    .io_data_2_out_valid(PE_256_io_data_2_out_valid),
    .io_data_2_out_bits(PE_256_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_256_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_256_io_data_1_in_valid),
    .io_data_1_in_bits(PE_256_io_data_1_in_bits),
    .io_data_1_out_valid(PE_256_io_data_1_out_valid),
    .io_data_1_out_bits(PE_256_io_data_1_out_bits),
    .io_data_0_in_valid(PE_256_io_data_0_in_valid),
    .io_data_0_in_bits(PE_256_io_data_0_in_bits),
    .io_data_0_out_valid(PE_256_io_data_0_out_valid),
    .io_data_0_out_bits(PE_256_io_data_0_out_bits)
  );
  PE PE_257 ( // @[pe.scala 187:13]
    .clock(PE_257_clock),
    .reset(PE_257_reset),
    .io_data_2_out_valid(PE_257_io_data_2_out_valid),
    .io_data_2_out_bits(PE_257_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_257_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_257_io_data_1_in_valid),
    .io_data_1_in_bits(PE_257_io_data_1_in_bits),
    .io_data_1_out_valid(PE_257_io_data_1_out_valid),
    .io_data_1_out_bits(PE_257_io_data_1_out_bits),
    .io_data_0_in_valid(PE_257_io_data_0_in_valid),
    .io_data_0_in_bits(PE_257_io_data_0_in_bits),
    .io_data_0_out_valid(PE_257_io_data_0_out_valid),
    .io_data_0_out_bits(PE_257_io_data_0_out_bits)
  );
  PE PE_258 ( // @[pe.scala 187:13]
    .clock(PE_258_clock),
    .reset(PE_258_reset),
    .io_data_2_out_valid(PE_258_io_data_2_out_valid),
    .io_data_2_out_bits(PE_258_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_258_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_258_io_data_1_in_valid),
    .io_data_1_in_bits(PE_258_io_data_1_in_bits),
    .io_data_1_out_valid(PE_258_io_data_1_out_valid),
    .io_data_1_out_bits(PE_258_io_data_1_out_bits),
    .io_data_0_in_valid(PE_258_io_data_0_in_valid),
    .io_data_0_in_bits(PE_258_io_data_0_in_bits),
    .io_data_0_out_valid(PE_258_io_data_0_out_valid),
    .io_data_0_out_bits(PE_258_io_data_0_out_bits)
  );
  PE PE_259 ( // @[pe.scala 187:13]
    .clock(PE_259_clock),
    .reset(PE_259_reset),
    .io_data_2_out_valid(PE_259_io_data_2_out_valid),
    .io_data_2_out_bits(PE_259_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_259_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_259_io_data_1_in_valid),
    .io_data_1_in_bits(PE_259_io_data_1_in_bits),
    .io_data_1_out_valid(PE_259_io_data_1_out_valid),
    .io_data_1_out_bits(PE_259_io_data_1_out_bits),
    .io_data_0_in_valid(PE_259_io_data_0_in_valid),
    .io_data_0_in_bits(PE_259_io_data_0_in_bits),
    .io_data_0_out_valid(PE_259_io_data_0_out_valid),
    .io_data_0_out_bits(PE_259_io_data_0_out_bits)
  );
  PE PE_260 ( // @[pe.scala 187:13]
    .clock(PE_260_clock),
    .reset(PE_260_reset),
    .io_data_2_out_valid(PE_260_io_data_2_out_valid),
    .io_data_2_out_bits(PE_260_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_260_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_260_io_data_1_in_valid),
    .io_data_1_in_bits(PE_260_io_data_1_in_bits),
    .io_data_1_out_valid(PE_260_io_data_1_out_valid),
    .io_data_1_out_bits(PE_260_io_data_1_out_bits),
    .io_data_0_in_valid(PE_260_io_data_0_in_valid),
    .io_data_0_in_bits(PE_260_io_data_0_in_bits),
    .io_data_0_out_valid(PE_260_io_data_0_out_valid),
    .io_data_0_out_bits(PE_260_io_data_0_out_bits)
  );
  PE PE_261 ( // @[pe.scala 187:13]
    .clock(PE_261_clock),
    .reset(PE_261_reset),
    .io_data_2_out_valid(PE_261_io_data_2_out_valid),
    .io_data_2_out_bits(PE_261_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_261_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_261_io_data_1_in_valid),
    .io_data_1_in_bits(PE_261_io_data_1_in_bits),
    .io_data_1_out_valid(PE_261_io_data_1_out_valid),
    .io_data_1_out_bits(PE_261_io_data_1_out_bits),
    .io_data_0_in_valid(PE_261_io_data_0_in_valid),
    .io_data_0_in_bits(PE_261_io_data_0_in_bits),
    .io_data_0_out_valid(PE_261_io_data_0_out_valid),
    .io_data_0_out_bits(PE_261_io_data_0_out_bits)
  );
  PE PE_262 ( // @[pe.scala 187:13]
    .clock(PE_262_clock),
    .reset(PE_262_reset),
    .io_data_2_out_valid(PE_262_io_data_2_out_valid),
    .io_data_2_out_bits(PE_262_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_262_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_262_io_data_1_in_valid),
    .io_data_1_in_bits(PE_262_io_data_1_in_bits),
    .io_data_1_out_valid(PE_262_io_data_1_out_valid),
    .io_data_1_out_bits(PE_262_io_data_1_out_bits),
    .io_data_0_in_valid(PE_262_io_data_0_in_valid),
    .io_data_0_in_bits(PE_262_io_data_0_in_bits),
    .io_data_0_out_valid(PE_262_io_data_0_out_valid),
    .io_data_0_out_bits(PE_262_io_data_0_out_bits)
  );
  PE PE_263 ( // @[pe.scala 187:13]
    .clock(PE_263_clock),
    .reset(PE_263_reset),
    .io_data_2_out_valid(PE_263_io_data_2_out_valid),
    .io_data_2_out_bits(PE_263_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_263_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_263_io_data_1_in_valid),
    .io_data_1_in_bits(PE_263_io_data_1_in_bits),
    .io_data_1_out_valid(PE_263_io_data_1_out_valid),
    .io_data_1_out_bits(PE_263_io_data_1_out_bits),
    .io_data_0_in_valid(PE_263_io_data_0_in_valid),
    .io_data_0_in_bits(PE_263_io_data_0_in_bits),
    .io_data_0_out_valid(PE_263_io_data_0_out_valid),
    .io_data_0_out_bits(PE_263_io_data_0_out_bits)
  );
  PE PE_264 ( // @[pe.scala 187:13]
    .clock(PE_264_clock),
    .reset(PE_264_reset),
    .io_data_2_out_valid(PE_264_io_data_2_out_valid),
    .io_data_2_out_bits(PE_264_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_264_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_264_io_data_1_in_valid),
    .io_data_1_in_bits(PE_264_io_data_1_in_bits),
    .io_data_1_out_valid(PE_264_io_data_1_out_valid),
    .io_data_1_out_bits(PE_264_io_data_1_out_bits),
    .io_data_0_in_valid(PE_264_io_data_0_in_valid),
    .io_data_0_in_bits(PE_264_io_data_0_in_bits),
    .io_data_0_out_valid(PE_264_io_data_0_out_valid),
    .io_data_0_out_bits(PE_264_io_data_0_out_bits)
  );
  PE PE_265 ( // @[pe.scala 187:13]
    .clock(PE_265_clock),
    .reset(PE_265_reset),
    .io_data_2_out_valid(PE_265_io_data_2_out_valid),
    .io_data_2_out_bits(PE_265_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_265_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_265_io_data_1_in_valid),
    .io_data_1_in_bits(PE_265_io_data_1_in_bits),
    .io_data_1_out_valid(PE_265_io_data_1_out_valid),
    .io_data_1_out_bits(PE_265_io_data_1_out_bits),
    .io_data_0_in_valid(PE_265_io_data_0_in_valid),
    .io_data_0_in_bits(PE_265_io_data_0_in_bits),
    .io_data_0_out_valid(PE_265_io_data_0_out_valid),
    .io_data_0_out_bits(PE_265_io_data_0_out_bits)
  );
  PE PE_266 ( // @[pe.scala 187:13]
    .clock(PE_266_clock),
    .reset(PE_266_reset),
    .io_data_2_out_valid(PE_266_io_data_2_out_valid),
    .io_data_2_out_bits(PE_266_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_266_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_266_io_data_1_in_valid),
    .io_data_1_in_bits(PE_266_io_data_1_in_bits),
    .io_data_1_out_valid(PE_266_io_data_1_out_valid),
    .io_data_1_out_bits(PE_266_io_data_1_out_bits),
    .io_data_0_in_valid(PE_266_io_data_0_in_valid),
    .io_data_0_in_bits(PE_266_io_data_0_in_bits),
    .io_data_0_out_valid(PE_266_io_data_0_out_valid),
    .io_data_0_out_bits(PE_266_io_data_0_out_bits)
  );
  PE PE_267 ( // @[pe.scala 187:13]
    .clock(PE_267_clock),
    .reset(PE_267_reset),
    .io_data_2_out_valid(PE_267_io_data_2_out_valid),
    .io_data_2_out_bits(PE_267_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_267_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_267_io_data_1_in_valid),
    .io_data_1_in_bits(PE_267_io_data_1_in_bits),
    .io_data_1_out_valid(PE_267_io_data_1_out_valid),
    .io_data_1_out_bits(PE_267_io_data_1_out_bits),
    .io_data_0_in_valid(PE_267_io_data_0_in_valid),
    .io_data_0_in_bits(PE_267_io_data_0_in_bits),
    .io_data_0_out_valid(PE_267_io_data_0_out_valid),
    .io_data_0_out_bits(PE_267_io_data_0_out_bits)
  );
  PE PE_268 ( // @[pe.scala 187:13]
    .clock(PE_268_clock),
    .reset(PE_268_reset),
    .io_data_2_out_valid(PE_268_io_data_2_out_valid),
    .io_data_2_out_bits(PE_268_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_268_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_268_io_data_1_in_valid),
    .io_data_1_in_bits(PE_268_io_data_1_in_bits),
    .io_data_1_out_valid(PE_268_io_data_1_out_valid),
    .io_data_1_out_bits(PE_268_io_data_1_out_bits),
    .io_data_0_in_valid(PE_268_io_data_0_in_valid),
    .io_data_0_in_bits(PE_268_io_data_0_in_bits),
    .io_data_0_out_valid(PE_268_io_data_0_out_valid),
    .io_data_0_out_bits(PE_268_io_data_0_out_bits)
  );
  PE PE_269 ( // @[pe.scala 187:13]
    .clock(PE_269_clock),
    .reset(PE_269_reset),
    .io_data_2_out_valid(PE_269_io_data_2_out_valid),
    .io_data_2_out_bits(PE_269_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_269_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_269_io_data_1_in_valid),
    .io_data_1_in_bits(PE_269_io_data_1_in_bits),
    .io_data_1_out_valid(PE_269_io_data_1_out_valid),
    .io_data_1_out_bits(PE_269_io_data_1_out_bits),
    .io_data_0_in_valid(PE_269_io_data_0_in_valid),
    .io_data_0_in_bits(PE_269_io_data_0_in_bits),
    .io_data_0_out_valid(PE_269_io_data_0_out_valid),
    .io_data_0_out_bits(PE_269_io_data_0_out_bits)
  );
  PE PE_270 ( // @[pe.scala 187:13]
    .clock(PE_270_clock),
    .reset(PE_270_reset),
    .io_data_2_out_valid(PE_270_io_data_2_out_valid),
    .io_data_2_out_bits(PE_270_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_270_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_270_io_data_1_in_valid),
    .io_data_1_in_bits(PE_270_io_data_1_in_bits),
    .io_data_1_out_valid(PE_270_io_data_1_out_valid),
    .io_data_1_out_bits(PE_270_io_data_1_out_bits),
    .io_data_0_in_valid(PE_270_io_data_0_in_valid),
    .io_data_0_in_bits(PE_270_io_data_0_in_bits),
    .io_data_0_out_valid(PE_270_io_data_0_out_valid),
    .io_data_0_out_bits(PE_270_io_data_0_out_bits)
  );
  PE PE_271 ( // @[pe.scala 187:13]
    .clock(PE_271_clock),
    .reset(PE_271_reset),
    .io_data_2_out_valid(PE_271_io_data_2_out_valid),
    .io_data_2_out_bits(PE_271_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_271_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_271_io_data_1_in_valid),
    .io_data_1_in_bits(PE_271_io_data_1_in_bits),
    .io_data_1_out_valid(PE_271_io_data_1_out_valid),
    .io_data_1_out_bits(PE_271_io_data_1_out_bits),
    .io_data_0_in_valid(PE_271_io_data_0_in_valid),
    .io_data_0_in_bits(PE_271_io_data_0_in_bits),
    .io_data_0_out_valid(PE_271_io_data_0_out_valid),
    .io_data_0_out_bits(PE_271_io_data_0_out_bits)
  );
  PE PE_272 ( // @[pe.scala 187:13]
    .clock(PE_272_clock),
    .reset(PE_272_reset),
    .io_data_2_out_valid(PE_272_io_data_2_out_valid),
    .io_data_2_out_bits(PE_272_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_272_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_272_io_data_1_in_valid),
    .io_data_1_in_bits(PE_272_io_data_1_in_bits),
    .io_data_1_out_valid(PE_272_io_data_1_out_valid),
    .io_data_1_out_bits(PE_272_io_data_1_out_bits),
    .io_data_0_in_valid(PE_272_io_data_0_in_valid),
    .io_data_0_in_bits(PE_272_io_data_0_in_bits),
    .io_data_0_out_valid(PE_272_io_data_0_out_valid),
    .io_data_0_out_bits(PE_272_io_data_0_out_bits)
  );
  PE PE_273 ( // @[pe.scala 187:13]
    .clock(PE_273_clock),
    .reset(PE_273_reset),
    .io_data_2_out_valid(PE_273_io_data_2_out_valid),
    .io_data_2_out_bits(PE_273_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_273_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_273_io_data_1_in_valid),
    .io_data_1_in_bits(PE_273_io_data_1_in_bits),
    .io_data_1_out_valid(PE_273_io_data_1_out_valid),
    .io_data_1_out_bits(PE_273_io_data_1_out_bits),
    .io_data_0_in_valid(PE_273_io_data_0_in_valid),
    .io_data_0_in_bits(PE_273_io_data_0_in_bits),
    .io_data_0_out_valid(PE_273_io_data_0_out_valid),
    .io_data_0_out_bits(PE_273_io_data_0_out_bits)
  );
  PE PE_274 ( // @[pe.scala 187:13]
    .clock(PE_274_clock),
    .reset(PE_274_reset),
    .io_data_2_out_valid(PE_274_io_data_2_out_valid),
    .io_data_2_out_bits(PE_274_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_274_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_274_io_data_1_in_valid),
    .io_data_1_in_bits(PE_274_io_data_1_in_bits),
    .io_data_1_out_valid(PE_274_io_data_1_out_valid),
    .io_data_1_out_bits(PE_274_io_data_1_out_bits),
    .io_data_0_in_valid(PE_274_io_data_0_in_valid),
    .io_data_0_in_bits(PE_274_io_data_0_in_bits),
    .io_data_0_out_valid(PE_274_io_data_0_out_valid),
    .io_data_0_out_bits(PE_274_io_data_0_out_bits)
  );
  PE PE_275 ( // @[pe.scala 187:13]
    .clock(PE_275_clock),
    .reset(PE_275_reset),
    .io_data_2_out_valid(PE_275_io_data_2_out_valid),
    .io_data_2_out_bits(PE_275_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_275_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_275_io_data_1_in_valid),
    .io_data_1_in_bits(PE_275_io_data_1_in_bits),
    .io_data_1_out_valid(PE_275_io_data_1_out_valid),
    .io_data_1_out_bits(PE_275_io_data_1_out_bits),
    .io_data_0_in_valid(PE_275_io_data_0_in_valid),
    .io_data_0_in_bits(PE_275_io_data_0_in_bits),
    .io_data_0_out_valid(PE_275_io_data_0_out_valid),
    .io_data_0_out_bits(PE_275_io_data_0_out_bits)
  );
  PE PE_276 ( // @[pe.scala 187:13]
    .clock(PE_276_clock),
    .reset(PE_276_reset),
    .io_data_2_out_valid(PE_276_io_data_2_out_valid),
    .io_data_2_out_bits(PE_276_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_276_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_276_io_data_1_in_valid),
    .io_data_1_in_bits(PE_276_io_data_1_in_bits),
    .io_data_1_out_valid(PE_276_io_data_1_out_valid),
    .io_data_1_out_bits(PE_276_io_data_1_out_bits),
    .io_data_0_in_valid(PE_276_io_data_0_in_valid),
    .io_data_0_in_bits(PE_276_io_data_0_in_bits),
    .io_data_0_out_valid(PE_276_io_data_0_out_valid),
    .io_data_0_out_bits(PE_276_io_data_0_out_bits)
  );
  PE PE_277 ( // @[pe.scala 187:13]
    .clock(PE_277_clock),
    .reset(PE_277_reset),
    .io_data_2_out_valid(PE_277_io_data_2_out_valid),
    .io_data_2_out_bits(PE_277_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_277_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_277_io_data_1_in_valid),
    .io_data_1_in_bits(PE_277_io_data_1_in_bits),
    .io_data_1_out_valid(PE_277_io_data_1_out_valid),
    .io_data_1_out_bits(PE_277_io_data_1_out_bits),
    .io_data_0_in_valid(PE_277_io_data_0_in_valid),
    .io_data_0_in_bits(PE_277_io_data_0_in_bits),
    .io_data_0_out_valid(PE_277_io_data_0_out_valid),
    .io_data_0_out_bits(PE_277_io_data_0_out_bits)
  );
  PE PE_278 ( // @[pe.scala 187:13]
    .clock(PE_278_clock),
    .reset(PE_278_reset),
    .io_data_2_out_valid(PE_278_io_data_2_out_valid),
    .io_data_2_out_bits(PE_278_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_278_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_278_io_data_1_in_valid),
    .io_data_1_in_bits(PE_278_io_data_1_in_bits),
    .io_data_1_out_valid(PE_278_io_data_1_out_valid),
    .io_data_1_out_bits(PE_278_io_data_1_out_bits),
    .io_data_0_in_valid(PE_278_io_data_0_in_valid),
    .io_data_0_in_bits(PE_278_io_data_0_in_bits),
    .io_data_0_out_valid(PE_278_io_data_0_out_valid),
    .io_data_0_out_bits(PE_278_io_data_0_out_bits)
  );
  PE PE_279 ( // @[pe.scala 187:13]
    .clock(PE_279_clock),
    .reset(PE_279_reset),
    .io_data_2_out_valid(PE_279_io_data_2_out_valid),
    .io_data_2_out_bits(PE_279_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_279_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_279_io_data_1_in_valid),
    .io_data_1_in_bits(PE_279_io_data_1_in_bits),
    .io_data_1_out_valid(PE_279_io_data_1_out_valid),
    .io_data_1_out_bits(PE_279_io_data_1_out_bits),
    .io_data_0_in_valid(PE_279_io_data_0_in_valid),
    .io_data_0_in_bits(PE_279_io_data_0_in_bits),
    .io_data_0_out_valid(PE_279_io_data_0_out_valid),
    .io_data_0_out_bits(PE_279_io_data_0_out_bits)
  );
  PE PE_280 ( // @[pe.scala 187:13]
    .clock(PE_280_clock),
    .reset(PE_280_reset),
    .io_data_2_out_valid(PE_280_io_data_2_out_valid),
    .io_data_2_out_bits(PE_280_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_280_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_280_io_data_1_in_valid),
    .io_data_1_in_bits(PE_280_io_data_1_in_bits),
    .io_data_1_out_valid(PE_280_io_data_1_out_valid),
    .io_data_1_out_bits(PE_280_io_data_1_out_bits),
    .io_data_0_in_valid(PE_280_io_data_0_in_valid),
    .io_data_0_in_bits(PE_280_io_data_0_in_bits),
    .io_data_0_out_valid(PE_280_io_data_0_out_valid),
    .io_data_0_out_bits(PE_280_io_data_0_out_bits)
  );
  PE PE_281 ( // @[pe.scala 187:13]
    .clock(PE_281_clock),
    .reset(PE_281_reset),
    .io_data_2_out_valid(PE_281_io_data_2_out_valid),
    .io_data_2_out_bits(PE_281_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_281_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_281_io_data_1_in_valid),
    .io_data_1_in_bits(PE_281_io_data_1_in_bits),
    .io_data_1_out_valid(PE_281_io_data_1_out_valid),
    .io_data_1_out_bits(PE_281_io_data_1_out_bits),
    .io_data_0_in_valid(PE_281_io_data_0_in_valid),
    .io_data_0_in_bits(PE_281_io_data_0_in_bits),
    .io_data_0_out_valid(PE_281_io_data_0_out_valid),
    .io_data_0_out_bits(PE_281_io_data_0_out_bits)
  );
  PE PE_282 ( // @[pe.scala 187:13]
    .clock(PE_282_clock),
    .reset(PE_282_reset),
    .io_data_2_out_valid(PE_282_io_data_2_out_valid),
    .io_data_2_out_bits(PE_282_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_282_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_282_io_data_1_in_valid),
    .io_data_1_in_bits(PE_282_io_data_1_in_bits),
    .io_data_1_out_valid(PE_282_io_data_1_out_valid),
    .io_data_1_out_bits(PE_282_io_data_1_out_bits),
    .io_data_0_in_valid(PE_282_io_data_0_in_valid),
    .io_data_0_in_bits(PE_282_io_data_0_in_bits),
    .io_data_0_out_valid(PE_282_io_data_0_out_valid),
    .io_data_0_out_bits(PE_282_io_data_0_out_bits)
  );
  PE PE_283 ( // @[pe.scala 187:13]
    .clock(PE_283_clock),
    .reset(PE_283_reset),
    .io_data_2_out_valid(PE_283_io_data_2_out_valid),
    .io_data_2_out_bits(PE_283_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_283_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_283_io_data_1_in_valid),
    .io_data_1_in_bits(PE_283_io_data_1_in_bits),
    .io_data_1_out_valid(PE_283_io_data_1_out_valid),
    .io_data_1_out_bits(PE_283_io_data_1_out_bits),
    .io_data_0_in_valid(PE_283_io_data_0_in_valid),
    .io_data_0_in_bits(PE_283_io_data_0_in_bits),
    .io_data_0_out_valid(PE_283_io_data_0_out_valid),
    .io_data_0_out_bits(PE_283_io_data_0_out_bits)
  );
  PE PE_284 ( // @[pe.scala 187:13]
    .clock(PE_284_clock),
    .reset(PE_284_reset),
    .io_data_2_out_valid(PE_284_io_data_2_out_valid),
    .io_data_2_out_bits(PE_284_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_284_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_284_io_data_1_in_valid),
    .io_data_1_in_bits(PE_284_io_data_1_in_bits),
    .io_data_1_out_valid(PE_284_io_data_1_out_valid),
    .io_data_1_out_bits(PE_284_io_data_1_out_bits),
    .io_data_0_in_valid(PE_284_io_data_0_in_valid),
    .io_data_0_in_bits(PE_284_io_data_0_in_bits),
    .io_data_0_out_valid(PE_284_io_data_0_out_valid),
    .io_data_0_out_bits(PE_284_io_data_0_out_bits)
  );
  PE PE_285 ( // @[pe.scala 187:13]
    .clock(PE_285_clock),
    .reset(PE_285_reset),
    .io_data_2_out_valid(PE_285_io_data_2_out_valid),
    .io_data_2_out_bits(PE_285_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_285_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_285_io_data_1_in_valid),
    .io_data_1_in_bits(PE_285_io_data_1_in_bits),
    .io_data_1_out_valid(PE_285_io_data_1_out_valid),
    .io_data_1_out_bits(PE_285_io_data_1_out_bits),
    .io_data_0_in_valid(PE_285_io_data_0_in_valid),
    .io_data_0_in_bits(PE_285_io_data_0_in_bits),
    .io_data_0_out_valid(PE_285_io_data_0_out_valid),
    .io_data_0_out_bits(PE_285_io_data_0_out_bits)
  );
  PE PE_286 ( // @[pe.scala 187:13]
    .clock(PE_286_clock),
    .reset(PE_286_reset),
    .io_data_2_out_valid(PE_286_io_data_2_out_valid),
    .io_data_2_out_bits(PE_286_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_286_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_286_io_data_1_in_valid),
    .io_data_1_in_bits(PE_286_io_data_1_in_bits),
    .io_data_1_out_valid(PE_286_io_data_1_out_valid),
    .io_data_1_out_bits(PE_286_io_data_1_out_bits),
    .io_data_0_in_valid(PE_286_io_data_0_in_valid),
    .io_data_0_in_bits(PE_286_io_data_0_in_bits),
    .io_data_0_out_valid(PE_286_io_data_0_out_valid),
    .io_data_0_out_bits(PE_286_io_data_0_out_bits)
  );
  PE PE_287 ( // @[pe.scala 187:13]
    .clock(PE_287_clock),
    .reset(PE_287_reset),
    .io_data_2_out_valid(PE_287_io_data_2_out_valid),
    .io_data_2_out_bits(PE_287_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_287_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_287_io_data_1_in_valid),
    .io_data_1_in_bits(PE_287_io_data_1_in_bits),
    .io_data_1_out_valid(PE_287_io_data_1_out_valid),
    .io_data_1_out_bits(PE_287_io_data_1_out_bits),
    .io_data_0_in_valid(PE_287_io_data_0_in_valid),
    .io_data_0_in_bits(PE_287_io_data_0_in_bits),
    .io_data_0_out_valid(PE_287_io_data_0_out_valid),
    .io_data_0_out_bits(PE_287_io_data_0_out_bits)
  );
  PE PE_288 ( // @[pe.scala 187:13]
    .clock(PE_288_clock),
    .reset(PE_288_reset),
    .io_data_2_out_valid(PE_288_io_data_2_out_valid),
    .io_data_2_out_bits(PE_288_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_288_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_288_io_data_1_in_valid),
    .io_data_1_in_bits(PE_288_io_data_1_in_bits),
    .io_data_1_out_valid(PE_288_io_data_1_out_valid),
    .io_data_1_out_bits(PE_288_io_data_1_out_bits),
    .io_data_0_in_valid(PE_288_io_data_0_in_valid),
    .io_data_0_in_bits(PE_288_io_data_0_in_bits),
    .io_data_0_out_valid(PE_288_io_data_0_out_valid),
    .io_data_0_out_bits(PE_288_io_data_0_out_bits)
  );
  PE PE_289 ( // @[pe.scala 187:13]
    .clock(PE_289_clock),
    .reset(PE_289_reset),
    .io_data_2_out_valid(PE_289_io_data_2_out_valid),
    .io_data_2_out_bits(PE_289_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_289_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_289_io_data_1_in_valid),
    .io_data_1_in_bits(PE_289_io_data_1_in_bits),
    .io_data_1_out_valid(PE_289_io_data_1_out_valid),
    .io_data_1_out_bits(PE_289_io_data_1_out_bits),
    .io_data_0_in_valid(PE_289_io_data_0_in_valid),
    .io_data_0_in_bits(PE_289_io_data_0_in_bits),
    .io_data_0_out_valid(PE_289_io_data_0_out_valid),
    .io_data_0_out_bits(PE_289_io_data_0_out_bits)
  );
  PE PE_290 ( // @[pe.scala 187:13]
    .clock(PE_290_clock),
    .reset(PE_290_reset),
    .io_data_2_out_valid(PE_290_io_data_2_out_valid),
    .io_data_2_out_bits(PE_290_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_290_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_290_io_data_1_in_valid),
    .io_data_1_in_bits(PE_290_io_data_1_in_bits),
    .io_data_1_out_valid(PE_290_io_data_1_out_valid),
    .io_data_1_out_bits(PE_290_io_data_1_out_bits),
    .io_data_0_in_valid(PE_290_io_data_0_in_valid),
    .io_data_0_in_bits(PE_290_io_data_0_in_bits),
    .io_data_0_out_valid(PE_290_io_data_0_out_valid),
    .io_data_0_out_bits(PE_290_io_data_0_out_bits)
  );
  PE PE_291 ( // @[pe.scala 187:13]
    .clock(PE_291_clock),
    .reset(PE_291_reset),
    .io_data_2_out_valid(PE_291_io_data_2_out_valid),
    .io_data_2_out_bits(PE_291_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_291_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_291_io_data_1_in_valid),
    .io_data_1_in_bits(PE_291_io_data_1_in_bits),
    .io_data_1_out_valid(PE_291_io_data_1_out_valid),
    .io_data_1_out_bits(PE_291_io_data_1_out_bits),
    .io_data_0_in_valid(PE_291_io_data_0_in_valid),
    .io_data_0_in_bits(PE_291_io_data_0_in_bits),
    .io_data_0_out_valid(PE_291_io_data_0_out_valid),
    .io_data_0_out_bits(PE_291_io_data_0_out_bits)
  );
  PE PE_292 ( // @[pe.scala 187:13]
    .clock(PE_292_clock),
    .reset(PE_292_reset),
    .io_data_2_out_valid(PE_292_io_data_2_out_valid),
    .io_data_2_out_bits(PE_292_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_292_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_292_io_data_1_in_valid),
    .io_data_1_in_bits(PE_292_io_data_1_in_bits),
    .io_data_1_out_valid(PE_292_io_data_1_out_valid),
    .io_data_1_out_bits(PE_292_io_data_1_out_bits),
    .io_data_0_in_valid(PE_292_io_data_0_in_valid),
    .io_data_0_in_bits(PE_292_io_data_0_in_bits),
    .io_data_0_out_valid(PE_292_io_data_0_out_valid),
    .io_data_0_out_bits(PE_292_io_data_0_out_bits)
  );
  PE PE_293 ( // @[pe.scala 187:13]
    .clock(PE_293_clock),
    .reset(PE_293_reset),
    .io_data_2_out_valid(PE_293_io_data_2_out_valid),
    .io_data_2_out_bits(PE_293_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_293_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_293_io_data_1_in_valid),
    .io_data_1_in_bits(PE_293_io_data_1_in_bits),
    .io_data_1_out_valid(PE_293_io_data_1_out_valid),
    .io_data_1_out_bits(PE_293_io_data_1_out_bits),
    .io_data_0_in_valid(PE_293_io_data_0_in_valid),
    .io_data_0_in_bits(PE_293_io_data_0_in_bits),
    .io_data_0_out_valid(PE_293_io_data_0_out_valid),
    .io_data_0_out_bits(PE_293_io_data_0_out_bits)
  );
  PE PE_294 ( // @[pe.scala 187:13]
    .clock(PE_294_clock),
    .reset(PE_294_reset),
    .io_data_2_out_valid(PE_294_io_data_2_out_valid),
    .io_data_2_out_bits(PE_294_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_294_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_294_io_data_1_in_valid),
    .io_data_1_in_bits(PE_294_io_data_1_in_bits),
    .io_data_1_out_valid(PE_294_io_data_1_out_valid),
    .io_data_1_out_bits(PE_294_io_data_1_out_bits),
    .io_data_0_in_valid(PE_294_io_data_0_in_valid),
    .io_data_0_in_bits(PE_294_io_data_0_in_bits),
    .io_data_0_out_valid(PE_294_io_data_0_out_valid),
    .io_data_0_out_bits(PE_294_io_data_0_out_bits)
  );
  PE PE_295 ( // @[pe.scala 187:13]
    .clock(PE_295_clock),
    .reset(PE_295_reset),
    .io_data_2_out_valid(PE_295_io_data_2_out_valid),
    .io_data_2_out_bits(PE_295_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_295_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_295_io_data_1_in_valid),
    .io_data_1_in_bits(PE_295_io_data_1_in_bits),
    .io_data_1_out_valid(PE_295_io_data_1_out_valid),
    .io_data_1_out_bits(PE_295_io_data_1_out_bits),
    .io_data_0_in_valid(PE_295_io_data_0_in_valid),
    .io_data_0_in_bits(PE_295_io_data_0_in_bits),
    .io_data_0_out_valid(PE_295_io_data_0_out_valid),
    .io_data_0_out_bits(PE_295_io_data_0_out_bits)
  );
  PE PE_296 ( // @[pe.scala 187:13]
    .clock(PE_296_clock),
    .reset(PE_296_reset),
    .io_data_2_out_valid(PE_296_io_data_2_out_valid),
    .io_data_2_out_bits(PE_296_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_296_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_296_io_data_1_in_valid),
    .io_data_1_in_bits(PE_296_io_data_1_in_bits),
    .io_data_1_out_valid(PE_296_io_data_1_out_valid),
    .io_data_1_out_bits(PE_296_io_data_1_out_bits),
    .io_data_0_in_valid(PE_296_io_data_0_in_valid),
    .io_data_0_in_bits(PE_296_io_data_0_in_bits),
    .io_data_0_out_valid(PE_296_io_data_0_out_valid),
    .io_data_0_out_bits(PE_296_io_data_0_out_bits)
  );
  PE PE_297 ( // @[pe.scala 187:13]
    .clock(PE_297_clock),
    .reset(PE_297_reset),
    .io_data_2_out_valid(PE_297_io_data_2_out_valid),
    .io_data_2_out_bits(PE_297_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_297_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_297_io_data_1_in_valid),
    .io_data_1_in_bits(PE_297_io_data_1_in_bits),
    .io_data_1_out_valid(PE_297_io_data_1_out_valid),
    .io_data_1_out_bits(PE_297_io_data_1_out_bits),
    .io_data_0_in_valid(PE_297_io_data_0_in_valid),
    .io_data_0_in_bits(PE_297_io_data_0_in_bits),
    .io_data_0_out_valid(PE_297_io_data_0_out_valid),
    .io_data_0_out_bits(PE_297_io_data_0_out_bits)
  );
  PE PE_298 ( // @[pe.scala 187:13]
    .clock(PE_298_clock),
    .reset(PE_298_reset),
    .io_data_2_out_valid(PE_298_io_data_2_out_valid),
    .io_data_2_out_bits(PE_298_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_298_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_298_io_data_1_in_valid),
    .io_data_1_in_bits(PE_298_io_data_1_in_bits),
    .io_data_1_out_valid(PE_298_io_data_1_out_valid),
    .io_data_1_out_bits(PE_298_io_data_1_out_bits),
    .io_data_0_in_valid(PE_298_io_data_0_in_valid),
    .io_data_0_in_bits(PE_298_io_data_0_in_bits),
    .io_data_0_out_valid(PE_298_io_data_0_out_valid),
    .io_data_0_out_bits(PE_298_io_data_0_out_bits)
  );
  PE PE_299 ( // @[pe.scala 187:13]
    .clock(PE_299_clock),
    .reset(PE_299_reset),
    .io_data_2_out_valid(PE_299_io_data_2_out_valid),
    .io_data_2_out_bits(PE_299_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_299_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_299_io_data_1_in_valid),
    .io_data_1_in_bits(PE_299_io_data_1_in_bits),
    .io_data_1_out_valid(PE_299_io_data_1_out_valid),
    .io_data_1_out_bits(PE_299_io_data_1_out_bits),
    .io_data_0_in_valid(PE_299_io_data_0_in_valid),
    .io_data_0_in_bits(PE_299_io_data_0_in_bits),
    .io_data_0_out_valid(PE_299_io_data_0_out_valid),
    .io_data_0_out_bits(PE_299_io_data_0_out_bits)
  );
  PE PE_300 ( // @[pe.scala 187:13]
    .clock(PE_300_clock),
    .reset(PE_300_reset),
    .io_data_2_out_valid(PE_300_io_data_2_out_valid),
    .io_data_2_out_bits(PE_300_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_300_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_300_io_data_1_in_valid),
    .io_data_1_in_bits(PE_300_io_data_1_in_bits),
    .io_data_1_out_valid(PE_300_io_data_1_out_valid),
    .io_data_1_out_bits(PE_300_io_data_1_out_bits),
    .io_data_0_in_valid(PE_300_io_data_0_in_valid),
    .io_data_0_in_bits(PE_300_io_data_0_in_bits),
    .io_data_0_out_valid(PE_300_io_data_0_out_valid),
    .io_data_0_out_bits(PE_300_io_data_0_out_bits)
  );
  PE PE_301 ( // @[pe.scala 187:13]
    .clock(PE_301_clock),
    .reset(PE_301_reset),
    .io_data_2_out_valid(PE_301_io_data_2_out_valid),
    .io_data_2_out_bits(PE_301_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_301_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_301_io_data_1_in_valid),
    .io_data_1_in_bits(PE_301_io_data_1_in_bits),
    .io_data_1_out_valid(PE_301_io_data_1_out_valid),
    .io_data_1_out_bits(PE_301_io_data_1_out_bits),
    .io_data_0_in_valid(PE_301_io_data_0_in_valid),
    .io_data_0_in_bits(PE_301_io_data_0_in_bits),
    .io_data_0_out_valid(PE_301_io_data_0_out_valid),
    .io_data_0_out_bits(PE_301_io_data_0_out_bits)
  );
  PE PE_302 ( // @[pe.scala 187:13]
    .clock(PE_302_clock),
    .reset(PE_302_reset),
    .io_data_2_out_valid(PE_302_io_data_2_out_valid),
    .io_data_2_out_bits(PE_302_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_302_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_302_io_data_1_in_valid),
    .io_data_1_in_bits(PE_302_io_data_1_in_bits),
    .io_data_1_out_valid(PE_302_io_data_1_out_valid),
    .io_data_1_out_bits(PE_302_io_data_1_out_bits),
    .io_data_0_in_valid(PE_302_io_data_0_in_valid),
    .io_data_0_in_bits(PE_302_io_data_0_in_bits),
    .io_data_0_out_valid(PE_302_io_data_0_out_valid),
    .io_data_0_out_bits(PE_302_io_data_0_out_bits)
  );
  PE PE_303 ( // @[pe.scala 187:13]
    .clock(PE_303_clock),
    .reset(PE_303_reset),
    .io_data_2_out_valid(PE_303_io_data_2_out_valid),
    .io_data_2_out_bits(PE_303_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_303_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_303_io_data_1_in_valid),
    .io_data_1_in_bits(PE_303_io_data_1_in_bits),
    .io_data_1_out_valid(PE_303_io_data_1_out_valid),
    .io_data_1_out_bits(PE_303_io_data_1_out_bits),
    .io_data_0_in_valid(PE_303_io_data_0_in_valid),
    .io_data_0_in_bits(PE_303_io_data_0_in_bits),
    .io_data_0_out_valid(PE_303_io_data_0_out_valid),
    .io_data_0_out_bits(PE_303_io_data_0_out_bits)
  );
  PE PE_304 ( // @[pe.scala 187:13]
    .clock(PE_304_clock),
    .reset(PE_304_reset),
    .io_data_2_out_valid(PE_304_io_data_2_out_valid),
    .io_data_2_out_bits(PE_304_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_304_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_304_io_data_1_in_valid),
    .io_data_1_in_bits(PE_304_io_data_1_in_bits),
    .io_data_1_out_valid(PE_304_io_data_1_out_valid),
    .io_data_1_out_bits(PE_304_io_data_1_out_bits),
    .io_data_0_in_valid(PE_304_io_data_0_in_valid),
    .io_data_0_in_bits(PE_304_io_data_0_in_bits),
    .io_data_0_out_valid(PE_304_io_data_0_out_valid),
    .io_data_0_out_bits(PE_304_io_data_0_out_bits)
  );
  PE PE_305 ( // @[pe.scala 187:13]
    .clock(PE_305_clock),
    .reset(PE_305_reset),
    .io_data_2_out_valid(PE_305_io_data_2_out_valid),
    .io_data_2_out_bits(PE_305_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_305_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_305_io_data_1_in_valid),
    .io_data_1_in_bits(PE_305_io_data_1_in_bits),
    .io_data_1_out_valid(PE_305_io_data_1_out_valid),
    .io_data_1_out_bits(PE_305_io_data_1_out_bits),
    .io_data_0_in_valid(PE_305_io_data_0_in_valid),
    .io_data_0_in_bits(PE_305_io_data_0_in_bits),
    .io_data_0_out_valid(PE_305_io_data_0_out_valid),
    .io_data_0_out_bits(PE_305_io_data_0_out_bits)
  );
  PE PE_306 ( // @[pe.scala 187:13]
    .clock(PE_306_clock),
    .reset(PE_306_reset),
    .io_data_2_out_valid(PE_306_io_data_2_out_valid),
    .io_data_2_out_bits(PE_306_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_306_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_306_io_data_1_in_valid),
    .io_data_1_in_bits(PE_306_io_data_1_in_bits),
    .io_data_1_out_valid(PE_306_io_data_1_out_valid),
    .io_data_1_out_bits(PE_306_io_data_1_out_bits),
    .io_data_0_in_valid(PE_306_io_data_0_in_valid),
    .io_data_0_in_bits(PE_306_io_data_0_in_bits),
    .io_data_0_out_valid(PE_306_io_data_0_out_valid),
    .io_data_0_out_bits(PE_306_io_data_0_out_bits)
  );
  PE PE_307 ( // @[pe.scala 187:13]
    .clock(PE_307_clock),
    .reset(PE_307_reset),
    .io_data_2_out_valid(PE_307_io_data_2_out_valid),
    .io_data_2_out_bits(PE_307_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_307_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_307_io_data_1_in_valid),
    .io_data_1_in_bits(PE_307_io_data_1_in_bits),
    .io_data_1_out_valid(PE_307_io_data_1_out_valid),
    .io_data_1_out_bits(PE_307_io_data_1_out_bits),
    .io_data_0_in_valid(PE_307_io_data_0_in_valid),
    .io_data_0_in_bits(PE_307_io_data_0_in_bits),
    .io_data_0_out_valid(PE_307_io_data_0_out_valid),
    .io_data_0_out_bits(PE_307_io_data_0_out_bits)
  );
  PE PE_308 ( // @[pe.scala 187:13]
    .clock(PE_308_clock),
    .reset(PE_308_reset),
    .io_data_2_out_valid(PE_308_io_data_2_out_valid),
    .io_data_2_out_bits(PE_308_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_308_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_308_io_data_1_in_valid),
    .io_data_1_in_bits(PE_308_io_data_1_in_bits),
    .io_data_1_out_valid(PE_308_io_data_1_out_valid),
    .io_data_1_out_bits(PE_308_io_data_1_out_bits),
    .io_data_0_in_valid(PE_308_io_data_0_in_valid),
    .io_data_0_in_bits(PE_308_io_data_0_in_bits),
    .io_data_0_out_valid(PE_308_io_data_0_out_valid),
    .io_data_0_out_bits(PE_308_io_data_0_out_bits)
  );
  PE PE_309 ( // @[pe.scala 187:13]
    .clock(PE_309_clock),
    .reset(PE_309_reset),
    .io_data_2_out_valid(PE_309_io_data_2_out_valid),
    .io_data_2_out_bits(PE_309_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_309_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_309_io_data_1_in_valid),
    .io_data_1_in_bits(PE_309_io_data_1_in_bits),
    .io_data_1_out_valid(PE_309_io_data_1_out_valid),
    .io_data_1_out_bits(PE_309_io_data_1_out_bits),
    .io_data_0_in_valid(PE_309_io_data_0_in_valid),
    .io_data_0_in_bits(PE_309_io_data_0_in_bits),
    .io_data_0_out_valid(PE_309_io_data_0_out_valid),
    .io_data_0_out_bits(PE_309_io_data_0_out_bits)
  );
  PE PE_310 ( // @[pe.scala 187:13]
    .clock(PE_310_clock),
    .reset(PE_310_reset),
    .io_data_2_out_valid(PE_310_io_data_2_out_valid),
    .io_data_2_out_bits(PE_310_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_310_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_310_io_data_1_in_valid),
    .io_data_1_in_bits(PE_310_io_data_1_in_bits),
    .io_data_1_out_valid(PE_310_io_data_1_out_valid),
    .io_data_1_out_bits(PE_310_io_data_1_out_bits),
    .io_data_0_in_valid(PE_310_io_data_0_in_valid),
    .io_data_0_in_bits(PE_310_io_data_0_in_bits),
    .io_data_0_out_valid(PE_310_io_data_0_out_valid),
    .io_data_0_out_bits(PE_310_io_data_0_out_bits)
  );
  PE PE_311 ( // @[pe.scala 187:13]
    .clock(PE_311_clock),
    .reset(PE_311_reset),
    .io_data_2_out_valid(PE_311_io_data_2_out_valid),
    .io_data_2_out_bits(PE_311_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_311_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_311_io_data_1_in_valid),
    .io_data_1_in_bits(PE_311_io_data_1_in_bits),
    .io_data_1_out_valid(PE_311_io_data_1_out_valid),
    .io_data_1_out_bits(PE_311_io_data_1_out_bits),
    .io_data_0_in_valid(PE_311_io_data_0_in_valid),
    .io_data_0_in_bits(PE_311_io_data_0_in_bits),
    .io_data_0_out_valid(PE_311_io_data_0_out_valid),
    .io_data_0_out_bits(PE_311_io_data_0_out_bits)
  );
  PE PE_312 ( // @[pe.scala 187:13]
    .clock(PE_312_clock),
    .reset(PE_312_reset),
    .io_data_2_out_valid(PE_312_io_data_2_out_valid),
    .io_data_2_out_bits(PE_312_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_312_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_312_io_data_1_in_valid),
    .io_data_1_in_bits(PE_312_io_data_1_in_bits),
    .io_data_1_out_valid(PE_312_io_data_1_out_valid),
    .io_data_1_out_bits(PE_312_io_data_1_out_bits),
    .io_data_0_in_valid(PE_312_io_data_0_in_valid),
    .io_data_0_in_bits(PE_312_io_data_0_in_bits),
    .io_data_0_out_valid(PE_312_io_data_0_out_valid),
    .io_data_0_out_bits(PE_312_io_data_0_out_bits)
  );
  PE PE_313 ( // @[pe.scala 187:13]
    .clock(PE_313_clock),
    .reset(PE_313_reset),
    .io_data_2_out_valid(PE_313_io_data_2_out_valid),
    .io_data_2_out_bits(PE_313_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_313_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_313_io_data_1_in_valid),
    .io_data_1_in_bits(PE_313_io_data_1_in_bits),
    .io_data_1_out_valid(PE_313_io_data_1_out_valid),
    .io_data_1_out_bits(PE_313_io_data_1_out_bits),
    .io_data_0_in_valid(PE_313_io_data_0_in_valid),
    .io_data_0_in_bits(PE_313_io_data_0_in_bits),
    .io_data_0_out_valid(PE_313_io_data_0_out_valid),
    .io_data_0_out_bits(PE_313_io_data_0_out_bits)
  );
  PE PE_314 ( // @[pe.scala 187:13]
    .clock(PE_314_clock),
    .reset(PE_314_reset),
    .io_data_2_out_valid(PE_314_io_data_2_out_valid),
    .io_data_2_out_bits(PE_314_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_314_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_314_io_data_1_in_valid),
    .io_data_1_in_bits(PE_314_io_data_1_in_bits),
    .io_data_1_out_valid(PE_314_io_data_1_out_valid),
    .io_data_1_out_bits(PE_314_io_data_1_out_bits),
    .io_data_0_in_valid(PE_314_io_data_0_in_valid),
    .io_data_0_in_bits(PE_314_io_data_0_in_bits),
    .io_data_0_out_valid(PE_314_io_data_0_out_valid),
    .io_data_0_out_bits(PE_314_io_data_0_out_bits)
  );
  PE PE_315 ( // @[pe.scala 187:13]
    .clock(PE_315_clock),
    .reset(PE_315_reset),
    .io_data_2_out_valid(PE_315_io_data_2_out_valid),
    .io_data_2_out_bits(PE_315_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_315_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_315_io_data_1_in_valid),
    .io_data_1_in_bits(PE_315_io_data_1_in_bits),
    .io_data_1_out_valid(PE_315_io_data_1_out_valid),
    .io_data_1_out_bits(PE_315_io_data_1_out_bits),
    .io_data_0_in_valid(PE_315_io_data_0_in_valid),
    .io_data_0_in_bits(PE_315_io_data_0_in_bits),
    .io_data_0_out_valid(PE_315_io_data_0_out_valid),
    .io_data_0_out_bits(PE_315_io_data_0_out_bits)
  );
  PE PE_316 ( // @[pe.scala 187:13]
    .clock(PE_316_clock),
    .reset(PE_316_reset),
    .io_data_2_out_valid(PE_316_io_data_2_out_valid),
    .io_data_2_out_bits(PE_316_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_316_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_316_io_data_1_in_valid),
    .io_data_1_in_bits(PE_316_io_data_1_in_bits),
    .io_data_1_out_valid(PE_316_io_data_1_out_valid),
    .io_data_1_out_bits(PE_316_io_data_1_out_bits),
    .io_data_0_in_valid(PE_316_io_data_0_in_valid),
    .io_data_0_in_bits(PE_316_io_data_0_in_bits),
    .io_data_0_out_valid(PE_316_io_data_0_out_valid),
    .io_data_0_out_bits(PE_316_io_data_0_out_bits)
  );
  PE PE_317 ( // @[pe.scala 187:13]
    .clock(PE_317_clock),
    .reset(PE_317_reset),
    .io_data_2_out_valid(PE_317_io_data_2_out_valid),
    .io_data_2_out_bits(PE_317_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_317_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_317_io_data_1_in_valid),
    .io_data_1_in_bits(PE_317_io_data_1_in_bits),
    .io_data_1_out_valid(PE_317_io_data_1_out_valid),
    .io_data_1_out_bits(PE_317_io_data_1_out_bits),
    .io_data_0_in_valid(PE_317_io_data_0_in_valid),
    .io_data_0_in_bits(PE_317_io_data_0_in_bits),
    .io_data_0_out_valid(PE_317_io_data_0_out_valid),
    .io_data_0_out_bits(PE_317_io_data_0_out_bits)
  );
  PE PE_318 ( // @[pe.scala 187:13]
    .clock(PE_318_clock),
    .reset(PE_318_reset),
    .io_data_2_out_valid(PE_318_io_data_2_out_valid),
    .io_data_2_out_bits(PE_318_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_318_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_318_io_data_1_in_valid),
    .io_data_1_in_bits(PE_318_io_data_1_in_bits),
    .io_data_1_out_valid(PE_318_io_data_1_out_valid),
    .io_data_1_out_bits(PE_318_io_data_1_out_bits),
    .io_data_0_in_valid(PE_318_io_data_0_in_valid),
    .io_data_0_in_bits(PE_318_io_data_0_in_bits),
    .io_data_0_out_valid(PE_318_io_data_0_out_valid),
    .io_data_0_out_bits(PE_318_io_data_0_out_bits)
  );
  PE PE_319 ( // @[pe.scala 187:13]
    .clock(PE_319_clock),
    .reset(PE_319_reset),
    .io_data_2_out_valid(PE_319_io_data_2_out_valid),
    .io_data_2_out_bits(PE_319_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_319_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_319_io_data_1_in_valid),
    .io_data_1_in_bits(PE_319_io_data_1_in_bits),
    .io_data_1_out_valid(PE_319_io_data_1_out_valid),
    .io_data_1_out_bits(PE_319_io_data_1_out_bits),
    .io_data_0_in_valid(PE_319_io_data_0_in_valid),
    .io_data_0_in_bits(PE_319_io_data_0_in_bits),
    .io_data_0_out_valid(PE_319_io_data_0_out_valid),
    .io_data_0_out_bits(PE_319_io_data_0_out_bits)
  );
  PE PE_320 ( // @[pe.scala 187:13]
    .clock(PE_320_clock),
    .reset(PE_320_reset),
    .io_data_2_out_valid(PE_320_io_data_2_out_valid),
    .io_data_2_out_bits(PE_320_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_320_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_320_io_data_1_in_valid),
    .io_data_1_in_bits(PE_320_io_data_1_in_bits),
    .io_data_1_out_valid(PE_320_io_data_1_out_valid),
    .io_data_1_out_bits(PE_320_io_data_1_out_bits),
    .io_data_0_in_valid(PE_320_io_data_0_in_valid),
    .io_data_0_in_bits(PE_320_io_data_0_in_bits),
    .io_data_0_out_valid(PE_320_io_data_0_out_valid),
    .io_data_0_out_bits(PE_320_io_data_0_out_bits)
  );
  PE PE_321 ( // @[pe.scala 187:13]
    .clock(PE_321_clock),
    .reset(PE_321_reset),
    .io_data_2_out_valid(PE_321_io_data_2_out_valid),
    .io_data_2_out_bits(PE_321_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_321_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_321_io_data_1_in_valid),
    .io_data_1_in_bits(PE_321_io_data_1_in_bits),
    .io_data_1_out_valid(PE_321_io_data_1_out_valid),
    .io_data_1_out_bits(PE_321_io_data_1_out_bits),
    .io_data_0_in_valid(PE_321_io_data_0_in_valid),
    .io_data_0_in_bits(PE_321_io_data_0_in_bits),
    .io_data_0_out_valid(PE_321_io_data_0_out_valid),
    .io_data_0_out_bits(PE_321_io_data_0_out_bits)
  );
  PE PE_322 ( // @[pe.scala 187:13]
    .clock(PE_322_clock),
    .reset(PE_322_reset),
    .io_data_2_out_valid(PE_322_io_data_2_out_valid),
    .io_data_2_out_bits(PE_322_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_322_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_322_io_data_1_in_valid),
    .io_data_1_in_bits(PE_322_io_data_1_in_bits),
    .io_data_1_out_valid(PE_322_io_data_1_out_valid),
    .io_data_1_out_bits(PE_322_io_data_1_out_bits),
    .io_data_0_in_valid(PE_322_io_data_0_in_valid),
    .io_data_0_in_bits(PE_322_io_data_0_in_bits),
    .io_data_0_out_valid(PE_322_io_data_0_out_valid),
    .io_data_0_out_bits(PE_322_io_data_0_out_bits)
  );
  PE PE_323 ( // @[pe.scala 187:13]
    .clock(PE_323_clock),
    .reset(PE_323_reset),
    .io_data_2_out_valid(PE_323_io_data_2_out_valid),
    .io_data_2_out_bits(PE_323_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_323_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_323_io_data_1_in_valid),
    .io_data_1_in_bits(PE_323_io_data_1_in_bits),
    .io_data_1_out_valid(PE_323_io_data_1_out_valid),
    .io_data_1_out_bits(PE_323_io_data_1_out_bits),
    .io_data_0_in_valid(PE_323_io_data_0_in_valid),
    .io_data_0_in_bits(PE_323_io_data_0_in_bits),
    .io_data_0_out_valid(PE_323_io_data_0_out_valid),
    .io_data_0_out_bits(PE_323_io_data_0_out_bits)
  );
  PE PE_324 ( // @[pe.scala 187:13]
    .clock(PE_324_clock),
    .reset(PE_324_reset),
    .io_data_2_out_valid(PE_324_io_data_2_out_valid),
    .io_data_2_out_bits(PE_324_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_324_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_324_io_data_1_in_valid),
    .io_data_1_in_bits(PE_324_io_data_1_in_bits),
    .io_data_1_out_valid(PE_324_io_data_1_out_valid),
    .io_data_1_out_bits(PE_324_io_data_1_out_bits),
    .io_data_0_in_valid(PE_324_io_data_0_in_valid),
    .io_data_0_in_bits(PE_324_io_data_0_in_bits),
    .io_data_0_out_valid(PE_324_io_data_0_out_valid),
    .io_data_0_out_bits(PE_324_io_data_0_out_bits)
  );
  PE PE_325 ( // @[pe.scala 187:13]
    .clock(PE_325_clock),
    .reset(PE_325_reset),
    .io_data_2_out_valid(PE_325_io_data_2_out_valid),
    .io_data_2_out_bits(PE_325_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_325_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_325_io_data_1_in_valid),
    .io_data_1_in_bits(PE_325_io_data_1_in_bits),
    .io_data_1_out_valid(PE_325_io_data_1_out_valid),
    .io_data_1_out_bits(PE_325_io_data_1_out_bits),
    .io_data_0_in_valid(PE_325_io_data_0_in_valid),
    .io_data_0_in_bits(PE_325_io_data_0_in_bits),
    .io_data_0_out_valid(PE_325_io_data_0_out_valid),
    .io_data_0_out_bits(PE_325_io_data_0_out_bits)
  );
  PE PE_326 ( // @[pe.scala 187:13]
    .clock(PE_326_clock),
    .reset(PE_326_reset),
    .io_data_2_out_valid(PE_326_io_data_2_out_valid),
    .io_data_2_out_bits(PE_326_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_326_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_326_io_data_1_in_valid),
    .io_data_1_in_bits(PE_326_io_data_1_in_bits),
    .io_data_1_out_valid(PE_326_io_data_1_out_valid),
    .io_data_1_out_bits(PE_326_io_data_1_out_bits),
    .io_data_0_in_valid(PE_326_io_data_0_in_valid),
    .io_data_0_in_bits(PE_326_io_data_0_in_bits),
    .io_data_0_out_valid(PE_326_io_data_0_out_valid),
    .io_data_0_out_bits(PE_326_io_data_0_out_bits)
  );
  PE PE_327 ( // @[pe.scala 187:13]
    .clock(PE_327_clock),
    .reset(PE_327_reset),
    .io_data_2_out_valid(PE_327_io_data_2_out_valid),
    .io_data_2_out_bits(PE_327_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_327_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_327_io_data_1_in_valid),
    .io_data_1_in_bits(PE_327_io_data_1_in_bits),
    .io_data_1_out_valid(PE_327_io_data_1_out_valid),
    .io_data_1_out_bits(PE_327_io_data_1_out_bits),
    .io_data_0_in_valid(PE_327_io_data_0_in_valid),
    .io_data_0_in_bits(PE_327_io_data_0_in_bits),
    .io_data_0_out_valid(PE_327_io_data_0_out_valid),
    .io_data_0_out_bits(PE_327_io_data_0_out_bits)
  );
  PE PE_328 ( // @[pe.scala 187:13]
    .clock(PE_328_clock),
    .reset(PE_328_reset),
    .io_data_2_out_valid(PE_328_io_data_2_out_valid),
    .io_data_2_out_bits(PE_328_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_328_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_328_io_data_1_in_valid),
    .io_data_1_in_bits(PE_328_io_data_1_in_bits),
    .io_data_1_out_valid(PE_328_io_data_1_out_valid),
    .io_data_1_out_bits(PE_328_io_data_1_out_bits),
    .io_data_0_in_valid(PE_328_io_data_0_in_valid),
    .io_data_0_in_bits(PE_328_io_data_0_in_bits),
    .io_data_0_out_valid(PE_328_io_data_0_out_valid),
    .io_data_0_out_bits(PE_328_io_data_0_out_bits)
  );
  PE PE_329 ( // @[pe.scala 187:13]
    .clock(PE_329_clock),
    .reset(PE_329_reset),
    .io_data_2_out_valid(PE_329_io_data_2_out_valid),
    .io_data_2_out_bits(PE_329_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_329_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_329_io_data_1_in_valid),
    .io_data_1_in_bits(PE_329_io_data_1_in_bits),
    .io_data_1_out_valid(PE_329_io_data_1_out_valid),
    .io_data_1_out_bits(PE_329_io_data_1_out_bits),
    .io_data_0_in_valid(PE_329_io_data_0_in_valid),
    .io_data_0_in_bits(PE_329_io_data_0_in_bits),
    .io_data_0_out_valid(PE_329_io_data_0_out_valid),
    .io_data_0_out_bits(PE_329_io_data_0_out_bits)
  );
  PE PE_330 ( // @[pe.scala 187:13]
    .clock(PE_330_clock),
    .reset(PE_330_reset),
    .io_data_2_out_valid(PE_330_io_data_2_out_valid),
    .io_data_2_out_bits(PE_330_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_330_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_330_io_data_1_in_valid),
    .io_data_1_in_bits(PE_330_io_data_1_in_bits),
    .io_data_1_out_valid(PE_330_io_data_1_out_valid),
    .io_data_1_out_bits(PE_330_io_data_1_out_bits),
    .io_data_0_in_valid(PE_330_io_data_0_in_valid),
    .io_data_0_in_bits(PE_330_io_data_0_in_bits),
    .io_data_0_out_valid(PE_330_io_data_0_out_valid),
    .io_data_0_out_bits(PE_330_io_data_0_out_bits)
  );
  PE PE_331 ( // @[pe.scala 187:13]
    .clock(PE_331_clock),
    .reset(PE_331_reset),
    .io_data_2_out_valid(PE_331_io_data_2_out_valid),
    .io_data_2_out_bits(PE_331_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_331_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_331_io_data_1_in_valid),
    .io_data_1_in_bits(PE_331_io_data_1_in_bits),
    .io_data_1_out_valid(PE_331_io_data_1_out_valid),
    .io_data_1_out_bits(PE_331_io_data_1_out_bits),
    .io_data_0_in_valid(PE_331_io_data_0_in_valid),
    .io_data_0_in_bits(PE_331_io_data_0_in_bits),
    .io_data_0_out_valid(PE_331_io_data_0_out_valid),
    .io_data_0_out_bits(PE_331_io_data_0_out_bits)
  );
  PE PE_332 ( // @[pe.scala 187:13]
    .clock(PE_332_clock),
    .reset(PE_332_reset),
    .io_data_2_out_valid(PE_332_io_data_2_out_valid),
    .io_data_2_out_bits(PE_332_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_332_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_332_io_data_1_in_valid),
    .io_data_1_in_bits(PE_332_io_data_1_in_bits),
    .io_data_1_out_valid(PE_332_io_data_1_out_valid),
    .io_data_1_out_bits(PE_332_io_data_1_out_bits),
    .io_data_0_in_valid(PE_332_io_data_0_in_valid),
    .io_data_0_in_bits(PE_332_io_data_0_in_bits),
    .io_data_0_out_valid(PE_332_io_data_0_out_valid),
    .io_data_0_out_bits(PE_332_io_data_0_out_bits)
  );
  PE PE_333 ( // @[pe.scala 187:13]
    .clock(PE_333_clock),
    .reset(PE_333_reset),
    .io_data_2_out_valid(PE_333_io_data_2_out_valid),
    .io_data_2_out_bits(PE_333_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_333_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_333_io_data_1_in_valid),
    .io_data_1_in_bits(PE_333_io_data_1_in_bits),
    .io_data_1_out_valid(PE_333_io_data_1_out_valid),
    .io_data_1_out_bits(PE_333_io_data_1_out_bits),
    .io_data_0_in_valid(PE_333_io_data_0_in_valid),
    .io_data_0_in_bits(PE_333_io_data_0_in_bits),
    .io_data_0_out_valid(PE_333_io_data_0_out_valid),
    .io_data_0_out_bits(PE_333_io_data_0_out_bits)
  );
  PE PE_334 ( // @[pe.scala 187:13]
    .clock(PE_334_clock),
    .reset(PE_334_reset),
    .io_data_2_out_valid(PE_334_io_data_2_out_valid),
    .io_data_2_out_bits(PE_334_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_334_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_334_io_data_1_in_valid),
    .io_data_1_in_bits(PE_334_io_data_1_in_bits),
    .io_data_1_out_valid(PE_334_io_data_1_out_valid),
    .io_data_1_out_bits(PE_334_io_data_1_out_bits),
    .io_data_0_in_valid(PE_334_io_data_0_in_valid),
    .io_data_0_in_bits(PE_334_io_data_0_in_bits),
    .io_data_0_out_valid(PE_334_io_data_0_out_valid),
    .io_data_0_out_bits(PE_334_io_data_0_out_bits)
  );
  PE PE_335 ( // @[pe.scala 187:13]
    .clock(PE_335_clock),
    .reset(PE_335_reset),
    .io_data_2_out_valid(PE_335_io_data_2_out_valid),
    .io_data_2_out_bits(PE_335_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_335_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_335_io_data_1_in_valid),
    .io_data_1_in_bits(PE_335_io_data_1_in_bits),
    .io_data_1_out_valid(PE_335_io_data_1_out_valid),
    .io_data_1_out_bits(PE_335_io_data_1_out_bits),
    .io_data_0_in_valid(PE_335_io_data_0_in_valid),
    .io_data_0_in_bits(PE_335_io_data_0_in_bits),
    .io_data_0_out_valid(PE_335_io_data_0_out_valid),
    .io_data_0_out_bits(PE_335_io_data_0_out_bits)
  );
  PE PE_336 ( // @[pe.scala 187:13]
    .clock(PE_336_clock),
    .reset(PE_336_reset),
    .io_data_2_out_valid(PE_336_io_data_2_out_valid),
    .io_data_2_out_bits(PE_336_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_336_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_336_io_data_1_in_valid),
    .io_data_1_in_bits(PE_336_io_data_1_in_bits),
    .io_data_1_out_valid(PE_336_io_data_1_out_valid),
    .io_data_1_out_bits(PE_336_io_data_1_out_bits),
    .io_data_0_in_valid(PE_336_io_data_0_in_valid),
    .io_data_0_in_bits(PE_336_io_data_0_in_bits),
    .io_data_0_out_valid(PE_336_io_data_0_out_valid),
    .io_data_0_out_bits(PE_336_io_data_0_out_bits)
  );
  PE PE_337 ( // @[pe.scala 187:13]
    .clock(PE_337_clock),
    .reset(PE_337_reset),
    .io_data_2_out_valid(PE_337_io_data_2_out_valid),
    .io_data_2_out_bits(PE_337_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_337_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_337_io_data_1_in_valid),
    .io_data_1_in_bits(PE_337_io_data_1_in_bits),
    .io_data_1_out_valid(PE_337_io_data_1_out_valid),
    .io_data_1_out_bits(PE_337_io_data_1_out_bits),
    .io_data_0_in_valid(PE_337_io_data_0_in_valid),
    .io_data_0_in_bits(PE_337_io_data_0_in_bits),
    .io_data_0_out_valid(PE_337_io_data_0_out_valid),
    .io_data_0_out_bits(PE_337_io_data_0_out_bits)
  );
  PE PE_338 ( // @[pe.scala 187:13]
    .clock(PE_338_clock),
    .reset(PE_338_reset),
    .io_data_2_out_valid(PE_338_io_data_2_out_valid),
    .io_data_2_out_bits(PE_338_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_338_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_338_io_data_1_in_valid),
    .io_data_1_in_bits(PE_338_io_data_1_in_bits),
    .io_data_1_out_valid(PE_338_io_data_1_out_valid),
    .io_data_1_out_bits(PE_338_io_data_1_out_bits),
    .io_data_0_in_valid(PE_338_io_data_0_in_valid),
    .io_data_0_in_bits(PE_338_io_data_0_in_bits),
    .io_data_0_out_valid(PE_338_io_data_0_out_valid),
    .io_data_0_out_bits(PE_338_io_data_0_out_bits)
  );
  PE PE_339 ( // @[pe.scala 187:13]
    .clock(PE_339_clock),
    .reset(PE_339_reset),
    .io_data_2_out_valid(PE_339_io_data_2_out_valid),
    .io_data_2_out_bits(PE_339_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_339_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_339_io_data_1_in_valid),
    .io_data_1_in_bits(PE_339_io_data_1_in_bits),
    .io_data_1_out_valid(PE_339_io_data_1_out_valid),
    .io_data_1_out_bits(PE_339_io_data_1_out_bits),
    .io_data_0_in_valid(PE_339_io_data_0_in_valid),
    .io_data_0_in_bits(PE_339_io_data_0_in_bits),
    .io_data_0_out_valid(PE_339_io_data_0_out_valid),
    .io_data_0_out_bits(PE_339_io_data_0_out_bits)
  );
  PE PE_340 ( // @[pe.scala 187:13]
    .clock(PE_340_clock),
    .reset(PE_340_reset),
    .io_data_2_out_valid(PE_340_io_data_2_out_valid),
    .io_data_2_out_bits(PE_340_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_340_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_340_io_data_1_in_valid),
    .io_data_1_in_bits(PE_340_io_data_1_in_bits),
    .io_data_1_out_valid(PE_340_io_data_1_out_valid),
    .io_data_1_out_bits(PE_340_io_data_1_out_bits),
    .io_data_0_in_valid(PE_340_io_data_0_in_valid),
    .io_data_0_in_bits(PE_340_io_data_0_in_bits),
    .io_data_0_out_valid(PE_340_io_data_0_out_valid),
    .io_data_0_out_bits(PE_340_io_data_0_out_bits)
  );
  PE PE_341 ( // @[pe.scala 187:13]
    .clock(PE_341_clock),
    .reset(PE_341_reset),
    .io_data_2_out_valid(PE_341_io_data_2_out_valid),
    .io_data_2_out_bits(PE_341_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_341_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_341_io_data_1_in_valid),
    .io_data_1_in_bits(PE_341_io_data_1_in_bits),
    .io_data_1_out_valid(PE_341_io_data_1_out_valid),
    .io_data_1_out_bits(PE_341_io_data_1_out_bits),
    .io_data_0_in_valid(PE_341_io_data_0_in_valid),
    .io_data_0_in_bits(PE_341_io_data_0_in_bits),
    .io_data_0_out_valid(PE_341_io_data_0_out_valid),
    .io_data_0_out_bits(PE_341_io_data_0_out_bits)
  );
  PE PE_342 ( // @[pe.scala 187:13]
    .clock(PE_342_clock),
    .reset(PE_342_reset),
    .io_data_2_out_valid(PE_342_io_data_2_out_valid),
    .io_data_2_out_bits(PE_342_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_342_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_342_io_data_1_in_valid),
    .io_data_1_in_bits(PE_342_io_data_1_in_bits),
    .io_data_1_out_valid(PE_342_io_data_1_out_valid),
    .io_data_1_out_bits(PE_342_io_data_1_out_bits),
    .io_data_0_in_valid(PE_342_io_data_0_in_valid),
    .io_data_0_in_bits(PE_342_io_data_0_in_bits),
    .io_data_0_out_valid(PE_342_io_data_0_out_valid),
    .io_data_0_out_bits(PE_342_io_data_0_out_bits)
  );
  PE PE_343 ( // @[pe.scala 187:13]
    .clock(PE_343_clock),
    .reset(PE_343_reset),
    .io_data_2_out_valid(PE_343_io_data_2_out_valid),
    .io_data_2_out_bits(PE_343_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_343_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_343_io_data_1_in_valid),
    .io_data_1_in_bits(PE_343_io_data_1_in_bits),
    .io_data_1_out_valid(PE_343_io_data_1_out_valid),
    .io_data_1_out_bits(PE_343_io_data_1_out_bits),
    .io_data_0_in_valid(PE_343_io_data_0_in_valid),
    .io_data_0_in_bits(PE_343_io_data_0_in_bits),
    .io_data_0_out_valid(PE_343_io_data_0_out_valid),
    .io_data_0_out_bits(PE_343_io_data_0_out_bits)
  );
  PE PE_344 ( // @[pe.scala 187:13]
    .clock(PE_344_clock),
    .reset(PE_344_reset),
    .io_data_2_out_valid(PE_344_io_data_2_out_valid),
    .io_data_2_out_bits(PE_344_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_344_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_344_io_data_1_in_valid),
    .io_data_1_in_bits(PE_344_io_data_1_in_bits),
    .io_data_1_out_valid(PE_344_io_data_1_out_valid),
    .io_data_1_out_bits(PE_344_io_data_1_out_bits),
    .io_data_0_in_valid(PE_344_io_data_0_in_valid),
    .io_data_0_in_bits(PE_344_io_data_0_in_bits),
    .io_data_0_out_valid(PE_344_io_data_0_out_valid),
    .io_data_0_out_bits(PE_344_io_data_0_out_bits)
  );
  PE PE_345 ( // @[pe.scala 187:13]
    .clock(PE_345_clock),
    .reset(PE_345_reset),
    .io_data_2_out_valid(PE_345_io_data_2_out_valid),
    .io_data_2_out_bits(PE_345_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_345_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_345_io_data_1_in_valid),
    .io_data_1_in_bits(PE_345_io_data_1_in_bits),
    .io_data_1_out_valid(PE_345_io_data_1_out_valid),
    .io_data_1_out_bits(PE_345_io_data_1_out_bits),
    .io_data_0_in_valid(PE_345_io_data_0_in_valid),
    .io_data_0_in_bits(PE_345_io_data_0_in_bits),
    .io_data_0_out_valid(PE_345_io_data_0_out_valid),
    .io_data_0_out_bits(PE_345_io_data_0_out_bits)
  );
  PE PE_346 ( // @[pe.scala 187:13]
    .clock(PE_346_clock),
    .reset(PE_346_reset),
    .io_data_2_out_valid(PE_346_io_data_2_out_valid),
    .io_data_2_out_bits(PE_346_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_346_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_346_io_data_1_in_valid),
    .io_data_1_in_bits(PE_346_io_data_1_in_bits),
    .io_data_1_out_valid(PE_346_io_data_1_out_valid),
    .io_data_1_out_bits(PE_346_io_data_1_out_bits),
    .io_data_0_in_valid(PE_346_io_data_0_in_valid),
    .io_data_0_in_bits(PE_346_io_data_0_in_bits),
    .io_data_0_out_valid(PE_346_io_data_0_out_valid),
    .io_data_0_out_bits(PE_346_io_data_0_out_bits)
  );
  PE PE_347 ( // @[pe.scala 187:13]
    .clock(PE_347_clock),
    .reset(PE_347_reset),
    .io_data_2_out_valid(PE_347_io_data_2_out_valid),
    .io_data_2_out_bits(PE_347_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_347_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_347_io_data_1_in_valid),
    .io_data_1_in_bits(PE_347_io_data_1_in_bits),
    .io_data_1_out_valid(PE_347_io_data_1_out_valid),
    .io_data_1_out_bits(PE_347_io_data_1_out_bits),
    .io_data_0_in_valid(PE_347_io_data_0_in_valid),
    .io_data_0_in_bits(PE_347_io_data_0_in_bits),
    .io_data_0_out_valid(PE_347_io_data_0_out_valid),
    .io_data_0_out_bits(PE_347_io_data_0_out_bits)
  );
  PE PE_348 ( // @[pe.scala 187:13]
    .clock(PE_348_clock),
    .reset(PE_348_reset),
    .io_data_2_out_valid(PE_348_io_data_2_out_valid),
    .io_data_2_out_bits(PE_348_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_348_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_348_io_data_1_in_valid),
    .io_data_1_in_bits(PE_348_io_data_1_in_bits),
    .io_data_1_out_valid(PE_348_io_data_1_out_valid),
    .io_data_1_out_bits(PE_348_io_data_1_out_bits),
    .io_data_0_in_valid(PE_348_io_data_0_in_valid),
    .io_data_0_in_bits(PE_348_io_data_0_in_bits),
    .io_data_0_out_valid(PE_348_io_data_0_out_valid),
    .io_data_0_out_bits(PE_348_io_data_0_out_bits)
  );
  PE PE_349 ( // @[pe.scala 187:13]
    .clock(PE_349_clock),
    .reset(PE_349_reset),
    .io_data_2_out_valid(PE_349_io_data_2_out_valid),
    .io_data_2_out_bits(PE_349_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_349_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_349_io_data_1_in_valid),
    .io_data_1_in_bits(PE_349_io_data_1_in_bits),
    .io_data_1_out_valid(PE_349_io_data_1_out_valid),
    .io_data_1_out_bits(PE_349_io_data_1_out_bits),
    .io_data_0_in_valid(PE_349_io_data_0_in_valid),
    .io_data_0_in_bits(PE_349_io_data_0_in_bits),
    .io_data_0_out_valid(PE_349_io_data_0_out_valid),
    .io_data_0_out_bits(PE_349_io_data_0_out_bits)
  );
  PE PE_350 ( // @[pe.scala 187:13]
    .clock(PE_350_clock),
    .reset(PE_350_reset),
    .io_data_2_out_valid(PE_350_io_data_2_out_valid),
    .io_data_2_out_bits(PE_350_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_350_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_350_io_data_1_in_valid),
    .io_data_1_in_bits(PE_350_io_data_1_in_bits),
    .io_data_1_out_valid(PE_350_io_data_1_out_valid),
    .io_data_1_out_bits(PE_350_io_data_1_out_bits),
    .io_data_0_in_valid(PE_350_io_data_0_in_valid),
    .io_data_0_in_bits(PE_350_io_data_0_in_bits),
    .io_data_0_out_valid(PE_350_io_data_0_out_valid),
    .io_data_0_out_bits(PE_350_io_data_0_out_bits)
  );
  PE PE_351 ( // @[pe.scala 187:13]
    .clock(PE_351_clock),
    .reset(PE_351_reset),
    .io_data_2_out_valid(PE_351_io_data_2_out_valid),
    .io_data_2_out_bits(PE_351_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_351_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_351_io_data_1_in_valid),
    .io_data_1_in_bits(PE_351_io_data_1_in_bits),
    .io_data_1_out_valid(PE_351_io_data_1_out_valid),
    .io_data_1_out_bits(PE_351_io_data_1_out_bits),
    .io_data_0_in_valid(PE_351_io_data_0_in_valid),
    .io_data_0_in_bits(PE_351_io_data_0_in_bits),
    .io_data_0_out_valid(PE_351_io_data_0_out_valid),
    .io_data_0_out_bits(PE_351_io_data_0_out_bits)
  );
  PE PE_352 ( // @[pe.scala 187:13]
    .clock(PE_352_clock),
    .reset(PE_352_reset),
    .io_data_2_out_valid(PE_352_io_data_2_out_valid),
    .io_data_2_out_bits(PE_352_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_352_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_352_io_data_1_in_valid),
    .io_data_1_in_bits(PE_352_io_data_1_in_bits),
    .io_data_1_out_valid(PE_352_io_data_1_out_valid),
    .io_data_1_out_bits(PE_352_io_data_1_out_bits),
    .io_data_0_in_valid(PE_352_io_data_0_in_valid),
    .io_data_0_in_bits(PE_352_io_data_0_in_bits),
    .io_data_0_out_valid(PE_352_io_data_0_out_valid),
    .io_data_0_out_bits(PE_352_io_data_0_out_bits)
  );
  PE PE_353 ( // @[pe.scala 187:13]
    .clock(PE_353_clock),
    .reset(PE_353_reset),
    .io_data_2_out_valid(PE_353_io_data_2_out_valid),
    .io_data_2_out_bits(PE_353_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_353_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_353_io_data_1_in_valid),
    .io_data_1_in_bits(PE_353_io_data_1_in_bits),
    .io_data_1_out_valid(PE_353_io_data_1_out_valid),
    .io_data_1_out_bits(PE_353_io_data_1_out_bits),
    .io_data_0_in_valid(PE_353_io_data_0_in_valid),
    .io_data_0_in_bits(PE_353_io_data_0_in_bits),
    .io_data_0_out_valid(PE_353_io_data_0_out_valid),
    .io_data_0_out_bits(PE_353_io_data_0_out_bits)
  );
  PE PE_354 ( // @[pe.scala 187:13]
    .clock(PE_354_clock),
    .reset(PE_354_reset),
    .io_data_2_out_valid(PE_354_io_data_2_out_valid),
    .io_data_2_out_bits(PE_354_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_354_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_354_io_data_1_in_valid),
    .io_data_1_in_bits(PE_354_io_data_1_in_bits),
    .io_data_1_out_valid(PE_354_io_data_1_out_valid),
    .io_data_1_out_bits(PE_354_io_data_1_out_bits),
    .io_data_0_in_valid(PE_354_io_data_0_in_valid),
    .io_data_0_in_bits(PE_354_io_data_0_in_bits),
    .io_data_0_out_valid(PE_354_io_data_0_out_valid),
    .io_data_0_out_bits(PE_354_io_data_0_out_bits)
  );
  PE PE_355 ( // @[pe.scala 187:13]
    .clock(PE_355_clock),
    .reset(PE_355_reset),
    .io_data_2_out_valid(PE_355_io_data_2_out_valid),
    .io_data_2_out_bits(PE_355_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_355_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_355_io_data_1_in_valid),
    .io_data_1_in_bits(PE_355_io_data_1_in_bits),
    .io_data_1_out_valid(PE_355_io_data_1_out_valid),
    .io_data_1_out_bits(PE_355_io_data_1_out_bits),
    .io_data_0_in_valid(PE_355_io_data_0_in_valid),
    .io_data_0_in_bits(PE_355_io_data_0_in_bits),
    .io_data_0_out_valid(PE_355_io_data_0_out_valid),
    .io_data_0_out_bits(PE_355_io_data_0_out_bits)
  );
  PE PE_356 ( // @[pe.scala 187:13]
    .clock(PE_356_clock),
    .reset(PE_356_reset),
    .io_data_2_out_valid(PE_356_io_data_2_out_valid),
    .io_data_2_out_bits(PE_356_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_356_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_356_io_data_1_in_valid),
    .io_data_1_in_bits(PE_356_io_data_1_in_bits),
    .io_data_1_out_valid(PE_356_io_data_1_out_valid),
    .io_data_1_out_bits(PE_356_io_data_1_out_bits),
    .io_data_0_in_valid(PE_356_io_data_0_in_valid),
    .io_data_0_in_bits(PE_356_io_data_0_in_bits),
    .io_data_0_out_valid(PE_356_io_data_0_out_valid),
    .io_data_0_out_bits(PE_356_io_data_0_out_bits)
  );
  PE PE_357 ( // @[pe.scala 187:13]
    .clock(PE_357_clock),
    .reset(PE_357_reset),
    .io_data_2_out_valid(PE_357_io_data_2_out_valid),
    .io_data_2_out_bits(PE_357_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_357_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_357_io_data_1_in_valid),
    .io_data_1_in_bits(PE_357_io_data_1_in_bits),
    .io_data_1_out_valid(PE_357_io_data_1_out_valid),
    .io_data_1_out_bits(PE_357_io_data_1_out_bits),
    .io_data_0_in_valid(PE_357_io_data_0_in_valid),
    .io_data_0_in_bits(PE_357_io_data_0_in_bits),
    .io_data_0_out_valid(PE_357_io_data_0_out_valid),
    .io_data_0_out_bits(PE_357_io_data_0_out_bits)
  );
  PE PE_358 ( // @[pe.scala 187:13]
    .clock(PE_358_clock),
    .reset(PE_358_reset),
    .io_data_2_out_valid(PE_358_io_data_2_out_valid),
    .io_data_2_out_bits(PE_358_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_358_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_358_io_data_1_in_valid),
    .io_data_1_in_bits(PE_358_io_data_1_in_bits),
    .io_data_1_out_valid(PE_358_io_data_1_out_valid),
    .io_data_1_out_bits(PE_358_io_data_1_out_bits),
    .io_data_0_in_valid(PE_358_io_data_0_in_valid),
    .io_data_0_in_bits(PE_358_io_data_0_in_bits),
    .io_data_0_out_valid(PE_358_io_data_0_out_valid),
    .io_data_0_out_bits(PE_358_io_data_0_out_bits)
  );
  PE PE_359 ( // @[pe.scala 187:13]
    .clock(PE_359_clock),
    .reset(PE_359_reset),
    .io_data_2_out_valid(PE_359_io_data_2_out_valid),
    .io_data_2_out_bits(PE_359_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_359_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_359_io_data_1_in_valid),
    .io_data_1_in_bits(PE_359_io_data_1_in_bits),
    .io_data_1_out_valid(PE_359_io_data_1_out_valid),
    .io_data_1_out_bits(PE_359_io_data_1_out_bits),
    .io_data_0_in_valid(PE_359_io_data_0_in_valid),
    .io_data_0_in_bits(PE_359_io_data_0_in_bits),
    .io_data_0_out_valid(PE_359_io_data_0_out_valid),
    .io_data_0_out_bits(PE_359_io_data_0_out_bits)
  );
  PE PE_360 ( // @[pe.scala 187:13]
    .clock(PE_360_clock),
    .reset(PE_360_reset),
    .io_data_2_out_valid(PE_360_io_data_2_out_valid),
    .io_data_2_out_bits(PE_360_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_360_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_360_io_data_1_in_valid),
    .io_data_1_in_bits(PE_360_io_data_1_in_bits),
    .io_data_1_out_valid(PE_360_io_data_1_out_valid),
    .io_data_1_out_bits(PE_360_io_data_1_out_bits),
    .io_data_0_in_valid(PE_360_io_data_0_in_valid),
    .io_data_0_in_bits(PE_360_io_data_0_in_bits),
    .io_data_0_out_valid(PE_360_io_data_0_out_valid),
    .io_data_0_out_bits(PE_360_io_data_0_out_bits)
  );
  PE PE_361 ( // @[pe.scala 187:13]
    .clock(PE_361_clock),
    .reset(PE_361_reset),
    .io_data_2_out_valid(PE_361_io_data_2_out_valid),
    .io_data_2_out_bits(PE_361_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_361_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_361_io_data_1_in_valid),
    .io_data_1_in_bits(PE_361_io_data_1_in_bits),
    .io_data_1_out_valid(PE_361_io_data_1_out_valid),
    .io_data_1_out_bits(PE_361_io_data_1_out_bits),
    .io_data_0_in_valid(PE_361_io_data_0_in_valid),
    .io_data_0_in_bits(PE_361_io_data_0_in_bits),
    .io_data_0_out_valid(PE_361_io_data_0_out_valid),
    .io_data_0_out_bits(PE_361_io_data_0_out_bits)
  );
  PE PE_362 ( // @[pe.scala 187:13]
    .clock(PE_362_clock),
    .reset(PE_362_reset),
    .io_data_2_out_valid(PE_362_io_data_2_out_valid),
    .io_data_2_out_bits(PE_362_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_362_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_362_io_data_1_in_valid),
    .io_data_1_in_bits(PE_362_io_data_1_in_bits),
    .io_data_1_out_valid(PE_362_io_data_1_out_valid),
    .io_data_1_out_bits(PE_362_io_data_1_out_bits),
    .io_data_0_in_valid(PE_362_io_data_0_in_valid),
    .io_data_0_in_bits(PE_362_io_data_0_in_bits),
    .io_data_0_out_valid(PE_362_io_data_0_out_valid),
    .io_data_0_out_bits(PE_362_io_data_0_out_bits)
  );
  PE PE_363 ( // @[pe.scala 187:13]
    .clock(PE_363_clock),
    .reset(PE_363_reset),
    .io_data_2_out_valid(PE_363_io_data_2_out_valid),
    .io_data_2_out_bits(PE_363_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_363_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_363_io_data_1_in_valid),
    .io_data_1_in_bits(PE_363_io_data_1_in_bits),
    .io_data_1_out_valid(PE_363_io_data_1_out_valid),
    .io_data_1_out_bits(PE_363_io_data_1_out_bits),
    .io_data_0_in_valid(PE_363_io_data_0_in_valid),
    .io_data_0_in_bits(PE_363_io_data_0_in_bits),
    .io_data_0_out_valid(PE_363_io_data_0_out_valid),
    .io_data_0_out_bits(PE_363_io_data_0_out_bits)
  );
  PE PE_364 ( // @[pe.scala 187:13]
    .clock(PE_364_clock),
    .reset(PE_364_reset),
    .io_data_2_out_valid(PE_364_io_data_2_out_valid),
    .io_data_2_out_bits(PE_364_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_364_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_364_io_data_1_in_valid),
    .io_data_1_in_bits(PE_364_io_data_1_in_bits),
    .io_data_1_out_valid(PE_364_io_data_1_out_valid),
    .io_data_1_out_bits(PE_364_io_data_1_out_bits),
    .io_data_0_in_valid(PE_364_io_data_0_in_valid),
    .io_data_0_in_bits(PE_364_io_data_0_in_bits),
    .io_data_0_out_valid(PE_364_io_data_0_out_valid),
    .io_data_0_out_bits(PE_364_io_data_0_out_bits)
  );
  PE PE_365 ( // @[pe.scala 187:13]
    .clock(PE_365_clock),
    .reset(PE_365_reset),
    .io_data_2_out_valid(PE_365_io_data_2_out_valid),
    .io_data_2_out_bits(PE_365_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_365_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_365_io_data_1_in_valid),
    .io_data_1_in_bits(PE_365_io_data_1_in_bits),
    .io_data_1_out_valid(PE_365_io_data_1_out_valid),
    .io_data_1_out_bits(PE_365_io_data_1_out_bits),
    .io_data_0_in_valid(PE_365_io_data_0_in_valid),
    .io_data_0_in_bits(PE_365_io_data_0_in_bits),
    .io_data_0_out_valid(PE_365_io_data_0_out_valid),
    .io_data_0_out_bits(PE_365_io_data_0_out_bits)
  );
  PE PE_366 ( // @[pe.scala 187:13]
    .clock(PE_366_clock),
    .reset(PE_366_reset),
    .io_data_2_out_valid(PE_366_io_data_2_out_valid),
    .io_data_2_out_bits(PE_366_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_366_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_366_io_data_1_in_valid),
    .io_data_1_in_bits(PE_366_io_data_1_in_bits),
    .io_data_1_out_valid(PE_366_io_data_1_out_valid),
    .io_data_1_out_bits(PE_366_io_data_1_out_bits),
    .io_data_0_in_valid(PE_366_io_data_0_in_valid),
    .io_data_0_in_bits(PE_366_io_data_0_in_bits),
    .io_data_0_out_valid(PE_366_io_data_0_out_valid),
    .io_data_0_out_bits(PE_366_io_data_0_out_bits)
  );
  PE PE_367 ( // @[pe.scala 187:13]
    .clock(PE_367_clock),
    .reset(PE_367_reset),
    .io_data_2_out_valid(PE_367_io_data_2_out_valid),
    .io_data_2_out_bits(PE_367_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_367_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_367_io_data_1_in_valid),
    .io_data_1_in_bits(PE_367_io_data_1_in_bits),
    .io_data_1_out_valid(PE_367_io_data_1_out_valid),
    .io_data_1_out_bits(PE_367_io_data_1_out_bits),
    .io_data_0_in_valid(PE_367_io_data_0_in_valid),
    .io_data_0_in_bits(PE_367_io_data_0_in_bits),
    .io_data_0_out_valid(PE_367_io_data_0_out_valid),
    .io_data_0_out_bits(PE_367_io_data_0_out_bits)
  );
  PE PE_368 ( // @[pe.scala 187:13]
    .clock(PE_368_clock),
    .reset(PE_368_reset),
    .io_data_2_out_valid(PE_368_io_data_2_out_valid),
    .io_data_2_out_bits(PE_368_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_368_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_368_io_data_1_in_valid),
    .io_data_1_in_bits(PE_368_io_data_1_in_bits),
    .io_data_1_out_valid(PE_368_io_data_1_out_valid),
    .io_data_1_out_bits(PE_368_io_data_1_out_bits),
    .io_data_0_in_valid(PE_368_io_data_0_in_valid),
    .io_data_0_in_bits(PE_368_io_data_0_in_bits),
    .io_data_0_out_valid(PE_368_io_data_0_out_valid),
    .io_data_0_out_bits(PE_368_io_data_0_out_bits)
  );
  PE PE_369 ( // @[pe.scala 187:13]
    .clock(PE_369_clock),
    .reset(PE_369_reset),
    .io_data_2_out_valid(PE_369_io_data_2_out_valid),
    .io_data_2_out_bits(PE_369_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_369_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_369_io_data_1_in_valid),
    .io_data_1_in_bits(PE_369_io_data_1_in_bits),
    .io_data_1_out_valid(PE_369_io_data_1_out_valid),
    .io_data_1_out_bits(PE_369_io_data_1_out_bits),
    .io_data_0_in_valid(PE_369_io_data_0_in_valid),
    .io_data_0_in_bits(PE_369_io_data_0_in_bits),
    .io_data_0_out_valid(PE_369_io_data_0_out_valid),
    .io_data_0_out_bits(PE_369_io_data_0_out_bits)
  );
  PE PE_370 ( // @[pe.scala 187:13]
    .clock(PE_370_clock),
    .reset(PE_370_reset),
    .io_data_2_out_valid(PE_370_io_data_2_out_valid),
    .io_data_2_out_bits(PE_370_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_370_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_370_io_data_1_in_valid),
    .io_data_1_in_bits(PE_370_io_data_1_in_bits),
    .io_data_1_out_valid(PE_370_io_data_1_out_valid),
    .io_data_1_out_bits(PE_370_io_data_1_out_bits),
    .io_data_0_in_valid(PE_370_io_data_0_in_valid),
    .io_data_0_in_bits(PE_370_io_data_0_in_bits),
    .io_data_0_out_valid(PE_370_io_data_0_out_valid),
    .io_data_0_out_bits(PE_370_io_data_0_out_bits)
  );
  PE PE_371 ( // @[pe.scala 187:13]
    .clock(PE_371_clock),
    .reset(PE_371_reset),
    .io_data_2_out_valid(PE_371_io_data_2_out_valid),
    .io_data_2_out_bits(PE_371_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_371_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_371_io_data_1_in_valid),
    .io_data_1_in_bits(PE_371_io_data_1_in_bits),
    .io_data_1_out_valid(PE_371_io_data_1_out_valid),
    .io_data_1_out_bits(PE_371_io_data_1_out_bits),
    .io_data_0_in_valid(PE_371_io_data_0_in_valid),
    .io_data_0_in_bits(PE_371_io_data_0_in_bits),
    .io_data_0_out_valid(PE_371_io_data_0_out_valid),
    .io_data_0_out_bits(PE_371_io_data_0_out_bits)
  );
  PE PE_372 ( // @[pe.scala 187:13]
    .clock(PE_372_clock),
    .reset(PE_372_reset),
    .io_data_2_out_valid(PE_372_io_data_2_out_valid),
    .io_data_2_out_bits(PE_372_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_372_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_372_io_data_1_in_valid),
    .io_data_1_in_bits(PE_372_io_data_1_in_bits),
    .io_data_1_out_valid(PE_372_io_data_1_out_valid),
    .io_data_1_out_bits(PE_372_io_data_1_out_bits),
    .io_data_0_in_valid(PE_372_io_data_0_in_valid),
    .io_data_0_in_bits(PE_372_io_data_0_in_bits),
    .io_data_0_out_valid(PE_372_io_data_0_out_valid),
    .io_data_0_out_bits(PE_372_io_data_0_out_bits)
  );
  PE PE_373 ( // @[pe.scala 187:13]
    .clock(PE_373_clock),
    .reset(PE_373_reset),
    .io_data_2_out_valid(PE_373_io_data_2_out_valid),
    .io_data_2_out_bits(PE_373_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_373_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_373_io_data_1_in_valid),
    .io_data_1_in_bits(PE_373_io_data_1_in_bits),
    .io_data_1_out_valid(PE_373_io_data_1_out_valid),
    .io_data_1_out_bits(PE_373_io_data_1_out_bits),
    .io_data_0_in_valid(PE_373_io_data_0_in_valid),
    .io_data_0_in_bits(PE_373_io_data_0_in_bits),
    .io_data_0_out_valid(PE_373_io_data_0_out_valid),
    .io_data_0_out_bits(PE_373_io_data_0_out_bits)
  );
  PE PE_374 ( // @[pe.scala 187:13]
    .clock(PE_374_clock),
    .reset(PE_374_reset),
    .io_data_2_out_valid(PE_374_io_data_2_out_valid),
    .io_data_2_out_bits(PE_374_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_374_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_374_io_data_1_in_valid),
    .io_data_1_in_bits(PE_374_io_data_1_in_bits),
    .io_data_1_out_valid(PE_374_io_data_1_out_valid),
    .io_data_1_out_bits(PE_374_io_data_1_out_bits),
    .io_data_0_in_valid(PE_374_io_data_0_in_valid),
    .io_data_0_in_bits(PE_374_io_data_0_in_bits),
    .io_data_0_out_valid(PE_374_io_data_0_out_valid),
    .io_data_0_out_bits(PE_374_io_data_0_out_bits)
  );
  PE PE_375 ( // @[pe.scala 187:13]
    .clock(PE_375_clock),
    .reset(PE_375_reset),
    .io_data_2_out_valid(PE_375_io_data_2_out_valid),
    .io_data_2_out_bits(PE_375_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_375_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_375_io_data_1_in_valid),
    .io_data_1_in_bits(PE_375_io_data_1_in_bits),
    .io_data_1_out_valid(PE_375_io_data_1_out_valid),
    .io_data_1_out_bits(PE_375_io_data_1_out_bits),
    .io_data_0_in_valid(PE_375_io_data_0_in_valid),
    .io_data_0_in_bits(PE_375_io_data_0_in_bits),
    .io_data_0_out_valid(PE_375_io_data_0_out_valid),
    .io_data_0_out_bits(PE_375_io_data_0_out_bits)
  );
  PE PE_376 ( // @[pe.scala 187:13]
    .clock(PE_376_clock),
    .reset(PE_376_reset),
    .io_data_2_out_valid(PE_376_io_data_2_out_valid),
    .io_data_2_out_bits(PE_376_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_376_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_376_io_data_1_in_valid),
    .io_data_1_in_bits(PE_376_io_data_1_in_bits),
    .io_data_1_out_valid(PE_376_io_data_1_out_valid),
    .io_data_1_out_bits(PE_376_io_data_1_out_bits),
    .io_data_0_in_valid(PE_376_io_data_0_in_valid),
    .io_data_0_in_bits(PE_376_io_data_0_in_bits),
    .io_data_0_out_valid(PE_376_io_data_0_out_valid),
    .io_data_0_out_bits(PE_376_io_data_0_out_bits)
  );
  PE PE_377 ( // @[pe.scala 187:13]
    .clock(PE_377_clock),
    .reset(PE_377_reset),
    .io_data_2_out_valid(PE_377_io_data_2_out_valid),
    .io_data_2_out_bits(PE_377_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_377_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_377_io_data_1_in_valid),
    .io_data_1_in_bits(PE_377_io_data_1_in_bits),
    .io_data_1_out_valid(PE_377_io_data_1_out_valid),
    .io_data_1_out_bits(PE_377_io_data_1_out_bits),
    .io_data_0_in_valid(PE_377_io_data_0_in_valid),
    .io_data_0_in_bits(PE_377_io_data_0_in_bits),
    .io_data_0_out_valid(PE_377_io_data_0_out_valid),
    .io_data_0_out_bits(PE_377_io_data_0_out_bits)
  );
  PE PE_378 ( // @[pe.scala 187:13]
    .clock(PE_378_clock),
    .reset(PE_378_reset),
    .io_data_2_out_valid(PE_378_io_data_2_out_valid),
    .io_data_2_out_bits(PE_378_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_378_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_378_io_data_1_in_valid),
    .io_data_1_in_bits(PE_378_io_data_1_in_bits),
    .io_data_1_out_valid(PE_378_io_data_1_out_valid),
    .io_data_1_out_bits(PE_378_io_data_1_out_bits),
    .io_data_0_in_valid(PE_378_io_data_0_in_valid),
    .io_data_0_in_bits(PE_378_io_data_0_in_bits),
    .io_data_0_out_valid(PE_378_io_data_0_out_valid),
    .io_data_0_out_bits(PE_378_io_data_0_out_bits)
  );
  PE PE_379 ( // @[pe.scala 187:13]
    .clock(PE_379_clock),
    .reset(PE_379_reset),
    .io_data_2_out_valid(PE_379_io_data_2_out_valid),
    .io_data_2_out_bits(PE_379_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_379_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_379_io_data_1_in_valid),
    .io_data_1_in_bits(PE_379_io_data_1_in_bits),
    .io_data_1_out_valid(PE_379_io_data_1_out_valid),
    .io_data_1_out_bits(PE_379_io_data_1_out_bits),
    .io_data_0_in_valid(PE_379_io_data_0_in_valid),
    .io_data_0_in_bits(PE_379_io_data_0_in_bits),
    .io_data_0_out_valid(PE_379_io_data_0_out_valid),
    .io_data_0_out_bits(PE_379_io_data_0_out_bits)
  );
  PE PE_380 ( // @[pe.scala 187:13]
    .clock(PE_380_clock),
    .reset(PE_380_reset),
    .io_data_2_out_valid(PE_380_io_data_2_out_valid),
    .io_data_2_out_bits(PE_380_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_380_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_380_io_data_1_in_valid),
    .io_data_1_in_bits(PE_380_io_data_1_in_bits),
    .io_data_1_out_valid(PE_380_io_data_1_out_valid),
    .io_data_1_out_bits(PE_380_io_data_1_out_bits),
    .io_data_0_in_valid(PE_380_io_data_0_in_valid),
    .io_data_0_in_bits(PE_380_io_data_0_in_bits),
    .io_data_0_out_valid(PE_380_io_data_0_out_valid),
    .io_data_0_out_bits(PE_380_io_data_0_out_bits)
  );
  PE PE_381 ( // @[pe.scala 187:13]
    .clock(PE_381_clock),
    .reset(PE_381_reset),
    .io_data_2_out_valid(PE_381_io_data_2_out_valid),
    .io_data_2_out_bits(PE_381_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_381_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_381_io_data_1_in_valid),
    .io_data_1_in_bits(PE_381_io_data_1_in_bits),
    .io_data_1_out_valid(PE_381_io_data_1_out_valid),
    .io_data_1_out_bits(PE_381_io_data_1_out_bits),
    .io_data_0_in_valid(PE_381_io_data_0_in_valid),
    .io_data_0_in_bits(PE_381_io_data_0_in_bits),
    .io_data_0_out_valid(PE_381_io_data_0_out_valid),
    .io_data_0_out_bits(PE_381_io_data_0_out_bits)
  );
  PE PE_382 ( // @[pe.scala 187:13]
    .clock(PE_382_clock),
    .reset(PE_382_reset),
    .io_data_2_out_valid(PE_382_io_data_2_out_valid),
    .io_data_2_out_bits(PE_382_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_382_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_382_io_data_1_in_valid),
    .io_data_1_in_bits(PE_382_io_data_1_in_bits),
    .io_data_1_out_valid(PE_382_io_data_1_out_valid),
    .io_data_1_out_bits(PE_382_io_data_1_out_bits),
    .io_data_0_in_valid(PE_382_io_data_0_in_valid),
    .io_data_0_in_bits(PE_382_io_data_0_in_bits),
    .io_data_0_out_valid(PE_382_io_data_0_out_valid),
    .io_data_0_out_bits(PE_382_io_data_0_out_bits)
  );
  PE PE_383 ( // @[pe.scala 187:13]
    .clock(PE_383_clock),
    .reset(PE_383_reset),
    .io_data_2_out_valid(PE_383_io_data_2_out_valid),
    .io_data_2_out_bits(PE_383_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_383_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_383_io_data_1_in_valid),
    .io_data_1_in_bits(PE_383_io_data_1_in_bits),
    .io_data_1_out_valid(PE_383_io_data_1_out_valid),
    .io_data_1_out_bits(PE_383_io_data_1_out_bits),
    .io_data_0_in_valid(PE_383_io_data_0_in_valid),
    .io_data_0_in_bits(PE_383_io_data_0_in_bits),
    .io_data_0_out_valid(PE_383_io_data_0_out_valid),
    .io_data_0_out_bits(PE_383_io_data_0_out_bits)
  );
  PE PE_384 ( // @[pe.scala 187:13]
    .clock(PE_384_clock),
    .reset(PE_384_reset),
    .io_data_2_out_valid(PE_384_io_data_2_out_valid),
    .io_data_2_out_bits(PE_384_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_384_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_384_io_data_1_in_valid),
    .io_data_1_in_bits(PE_384_io_data_1_in_bits),
    .io_data_1_out_valid(PE_384_io_data_1_out_valid),
    .io_data_1_out_bits(PE_384_io_data_1_out_bits),
    .io_data_0_in_valid(PE_384_io_data_0_in_valid),
    .io_data_0_in_bits(PE_384_io_data_0_in_bits),
    .io_data_0_out_valid(PE_384_io_data_0_out_valid),
    .io_data_0_out_bits(PE_384_io_data_0_out_bits)
  );
  PE PE_385 ( // @[pe.scala 187:13]
    .clock(PE_385_clock),
    .reset(PE_385_reset),
    .io_data_2_out_valid(PE_385_io_data_2_out_valid),
    .io_data_2_out_bits(PE_385_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_385_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_385_io_data_1_in_valid),
    .io_data_1_in_bits(PE_385_io_data_1_in_bits),
    .io_data_1_out_valid(PE_385_io_data_1_out_valid),
    .io_data_1_out_bits(PE_385_io_data_1_out_bits),
    .io_data_0_in_valid(PE_385_io_data_0_in_valid),
    .io_data_0_in_bits(PE_385_io_data_0_in_bits),
    .io_data_0_out_valid(PE_385_io_data_0_out_valid),
    .io_data_0_out_bits(PE_385_io_data_0_out_bits)
  );
  PE PE_386 ( // @[pe.scala 187:13]
    .clock(PE_386_clock),
    .reset(PE_386_reset),
    .io_data_2_out_valid(PE_386_io_data_2_out_valid),
    .io_data_2_out_bits(PE_386_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_386_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_386_io_data_1_in_valid),
    .io_data_1_in_bits(PE_386_io_data_1_in_bits),
    .io_data_1_out_valid(PE_386_io_data_1_out_valid),
    .io_data_1_out_bits(PE_386_io_data_1_out_bits),
    .io_data_0_in_valid(PE_386_io_data_0_in_valid),
    .io_data_0_in_bits(PE_386_io_data_0_in_bits),
    .io_data_0_out_valid(PE_386_io_data_0_out_valid),
    .io_data_0_out_bits(PE_386_io_data_0_out_bits)
  );
  PE PE_387 ( // @[pe.scala 187:13]
    .clock(PE_387_clock),
    .reset(PE_387_reset),
    .io_data_2_out_valid(PE_387_io_data_2_out_valid),
    .io_data_2_out_bits(PE_387_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_387_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_387_io_data_1_in_valid),
    .io_data_1_in_bits(PE_387_io_data_1_in_bits),
    .io_data_1_out_valid(PE_387_io_data_1_out_valid),
    .io_data_1_out_bits(PE_387_io_data_1_out_bits),
    .io_data_0_in_valid(PE_387_io_data_0_in_valid),
    .io_data_0_in_bits(PE_387_io_data_0_in_bits),
    .io_data_0_out_valid(PE_387_io_data_0_out_valid),
    .io_data_0_out_bits(PE_387_io_data_0_out_bits)
  );
  PE PE_388 ( // @[pe.scala 187:13]
    .clock(PE_388_clock),
    .reset(PE_388_reset),
    .io_data_2_out_valid(PE_388_io_data_2_out_valid),
    .io_data_2_out_bits(PE_388_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_388_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_388_io_data_1_in_valid),
    .io_data_1_in_bits(PE_388_io_data_1_in_bits),
    .io_data_1_out_valid(PE_388_io_data_1_out_valid),
    .io_data_1_out_bits(PE_388_io_data_1_out_bits),
    .io_data_0_in_valid(PE_388_io_data_0_in_valid),
    .io_data_0_in_bits(PE_388_io_data_0_in_bits),
    .io_data_0_out_valid(PE_388_io_data_0_out_valid),
    .io_data_0_out_bits(PE_388_io_data_0_out_bits)
  );
  PE PE_389 ( // @[pe.scala 187:13]
    .clock(PE_389_clock),
    .reset(PE_389_reset),
    .io_data_2_out_valid(PE_389_io_data_2_out_valid),
    .io_data_2_out_bits(PE_389_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_389_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_389_io_data_1_in_valid),
    .io_data_1_in_bits(PE_389_io_data_1_in_bits),
    .io_data_1_out_valid(PE_389_io_data_1_out_valid),
    .io_data_1_out_bits(PE_389_io_data_1_out_bits),
    .io_data_0_in_valid(PE_389_io_data_0_in_valid),
    .io_data_0_in_bits(PE_389_io_data_0_in_bits),
    .io_data_0_out_valid(PE_389_io_data_0_out_valid),
    .io_data_0_out_bits(PE_389_io_data_0_out_bits)
  );
  PE PE_390 ( // @[pe.scala 187:13]
    .clock(PE_390_clock),
    .reset(PE_390_reset),
    .io_data_2_out_valid(PE_390_io_data_2_out_valid),
    .io_data_2_out_bits(PE_390_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_390_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_390_io_data_1_in_valid),
    .io_data_1_in_bits(PE_390_io_data_1_in_bits),
    .io_data_1_out_valid(PE_390_io_data_1_out_valid),
    .io_data_1_out_bits(PE_390_io_data_1_out_bits),
    .io_data_0_in_valid(PE_390_io_data_0_in_valid),
    .io_data_0_in_bits(PE_390_io_data_0_in_bits),
    .io_data_0_out_valid(PE_390_io_data_0_out_valid),
    .io_data_0_out_bits(PE_390_io_data_0_out_bits)
  );
  PE PE_391 ( // @[pe.scala 187:13]
    .clock(PE_391_clock),
    .reset(PE_391_reset),
    .io_data_2_out_valid(PE_391_io_data_2_out_valid),
    .io_data_2_out_bits(PE_391_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_391_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_391_io_data_1_in_valid),
    .io_data_1_in_bits(PE_391_io_data_1_in_bits),
    .io_data_1_out_valid(PE_391_io_data_1_out_valid),
    .io_data_1_out_bits(PE_391_io_data_1_out_bits),
    .io_data_0_in_valid(PE_391_io_data_0_in_valid),
    .io_data_0_in_bits(PE_391_io_data_0_in_bits),
    .io_data_0_out_valid(PE_391_io_data_0_out_valid),
    .io_data_0_out_bits(PE_391_io_data_0_out_bits)
  );
  PE PE_392 ( // @[pe.scala 187:13]
    .clock(PE_392_clock),
    .reset(PE_392_reset),
    .io_data_2_out_valid(PE_392_io_data_2_out_valid),
    .io_data_2_out_bits(PE_392_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_392_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_392_io_data_1_in_valid),
    .io_data_1_in_bits(PE_392_io_data_1_in_bits),
    .io_data_1_out_valid(PE_392_io_data_1_out_valid),
    .io_data_1_out_bits(PE_392_io_data_1_out_bits),
    .io_data_0_in_valid(PE_392_io_data_0_in_valid),
    .io_data_0_in_bits(PE_392_io_data_0_in_bits),
    .io_data_0_out_valid(PE_392_io_data_0_out_valid),
    .io_data_0_out_bits(PE_392_io_data_0_out_bits)
  );
  PE PE_393 ( // @[pe.scala 187:13]
    .clock(PE_393_clock),
    .reset(PE_393_reset),
    .io_data_2_out_valid(PE_393_io_data_2_out_valid),
    .io_data_2_out_bits(PE_393_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_393_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_393_io_data_1_in_valid),
    .io_data_1_in_bits(PE_393_io_data_1_in_bits),
    .io_data_1_out_valid(PE_393_io_data_1_out_valid),
    .io_data_1_out_bits(PE_393_io_data_1_out_bits),
    .io_data_0_in_valid(PE_393_io_data_0_in_valid),
    .io_data_0_in_bits(PE_393_io_data_0_in_bits),
    .io_data_0_out_valid(PE_393_io_data_0_out_valid),
    .io_data_0_out_bits(PE_393_io_data_0_out_bits)
  );
  PE PE_394 ( // @[pe.scala 187:13]
    .clock(PE_394_clock),
    .reset(PE_394_reset),
    .io_data_2_out_valid(PE_394_io_data_2_out_valid),
    .io_data_2_out_bits(PE_394_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_394_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_394_io_data_1_in_valid),
    .io_data_1_in_bits(PE_394_io_data_1_in_bits),
    .io_data_1_out_valid(PE_394_io_data_1_out_valid),
    .io_data_1_out_bits(PE_394_io_data_1_out_bits),
    .io_data_0_in_valid(PE_394_io_data_0_in_valid),
    .io_data_0_in_bits(PE_394_io_data_0_in_bits),
    .io_data_0_out_valid(PE_394_io_data_0_out_valid),
    .io_data_0_out_bits(PE_394_io_data_0_out_bits)
  );
  PE PE_395 ( // @[pe.scala 187:13]
    .clock(PE_395_clock),
    .reset(PE_395_reset),
    .io_data_2_out_valid(PE_395_io_data_2_out_valid),
    .io_data_2_out_bits(PE_395_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_395_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_395_io_data_1_in_valid),
    .io_data_1_in_bits(PE_395_io_data_1_in_bits),
    .io_data_1_out_valid(PE_395_io_data_1_out_valid),
    .io_data_1_out_bits(PE_395_io_data_1_out_bits),
    .io_data_0_in_valid(PE_395_io_data_0_in_valid),
    .io_data_0_in_bits(PE_395_io_data_0_in_bits),
    .io_data_0_out_valid(PE_395_io_data_0_out_valid),
    .io_data_0_out_bits(PE_395_io_data_0_out_bits)
  );
  PE PE_396 ( // @[pe.scala 187:13]
    .clock(PE_396_clock),
    .reset(PE_396_reset),
    .io_data_2_out_valid(PE_396_io_data_2_out_valid),
    .io_data_2_out_bits(PE_396_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_396_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_396_io_data_1_in_valid),
    .io_data_1_in_bits(PE_396_io_data_1_in_bits),
    .io_data_1_out_valid(PE_396_io_data_1_out_valid),
    .io_data_1_out_bits(PE_396_io_data_1_out_bits),
    .io_data_0_in_valid(PE_396_io_data_0_in_valid),
    .io_data_0_in_bits(PE_396_io_data_0_in_bits),
    .io_data_0_out_valid(PE_396_io_data_0_out_valid),
    .io_data_0_out_bits(PE_396_io_data_0_out_bits)
  );
  PE PE_397 ( // @[pe.scala 187:13]
    .clock(PE_397_clock),
    .reset(PE_397_reset),
    .io_data_2_out_valid(PE_397_io_data_2_out_valid),
    .io_data_2_out_bits(PE_397_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_397_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_397_io_data_1_in_valid),
    .io_data_1_in_bits(PE_397_io_data_1_in_bits),
    .io_data_1_out_valid(PE_397_io_data_1_out_valid),
    .io_data_1_out_bits(PE_397_io_data_1_out_bits),
    .io_data_0_in_valid(PE_397_io_data_0_in_valid),
    .io_data_0_in_bits(PE_397_io_data_0_in_bits),
    .io_data_0_out_valid(PE_397_io_data_0_out_valid),
    .io_data_0_out_bits(PE_397_io_data_0_out_bits)
  );
  PE PE_398 ( // @[pe.scala 187:13]
    .clock(PE_398_clock),
    .reset(PE_398_reset),
    .io_data_2_out_valid(PE_398_io_data_2_out_valid),
    .io_data_2_out_bits(PE_398_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_398_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_398_io_data_1_in_valid),
    .io_data_1_in_bits(PE_398_io_data_1_in_bits),
    .io_data_1_out_valid(PE_398_io_data_1_out_valid),
    .io_data_1_out_bits(PE_398_io_data_1_out_bits),
    .io_data_0_in_valid(PE_398_io_data_0_in_valid),
    .io_data_0_in_bits(PE_398_io_data_0_in_bits),
    .io_data_0_out_valid(PE_398_io_data_0_out_valid),
    .io_data_0_out_bits(PE_398_io_data_0_out_bits)
  );
  PE PE_399 ( // @[pe.scala 187:13]
    .clock(PE_399_clock),
    .reset(PE_399_reset),
    .io_data_2_out_valid(PE_399_io_data_2_out_valid),
    .io_data_2_out_bits(PE_399_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_399_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_399_io_data_1_in_valid),
    .io_data_1_in_bits(PE_399_io_data_1_in_bits),
    .io_data_1_out_valid(PE_399_io_data_1_out_valid),
    .io_data_1_out_bits(PE_399_io_data_1_out_bits),
    .io_data_0_in_valid(PE_399_io_data_0_in_valid),
    .io_data_0_in_bits(PE_399_io_data_0_in_bits),
    .io_data_0_out_valid(PE_399_io_data_0_out_valid),
    .io_data_0_out_bits(PE_399_io_data_0_out_bits)
  );
  PE PE_400 ( // @[pe.scala 187:13]
    .clock(PE_400_clock),
    .reset(PE_400_reset),
    .io_data_2_out_valid(PE_400_io_data_2_out_valid),
    .io_data_2_out_bits(PE_400_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_400_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_400_io_data_1_in_valid),
    .io_data_1_in_bits(PE_400_io_data_1_in_bits),
    .io_data_1_out_valid(PE_400_io_data_1_out_valid),
    .io_data_1_out_bits(PE_400_io_data_1_out_bits),
    .io_data_0_in_valid(PE_400_io_data_0_in_valid),
    .io_data_0_in_bits(PE_400_io_data_0_in_bits),
    .io_data_0_out_valid(PE_400_io_data_0_out_valid),
    .io_data_0_out_bits(PE_400_io_data_0_out_bits)
  );
  PE PE_401 ( // @[pe.scala 187:13]
    .clock(PE_401_clock),
    .reset(PE_401_reset),
    .io_data_2_out_valid(PE_401_io_data_2_out_valid),
    .io_data_2_out_bits(PE_401_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_401_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_401_io_data_1_in_valid),
    .io_data_1_in_bits(PE_401_io_data_1_in_bits),
    .io_data_1_out_valid(PE_401_io_data_1_out_valid),
    .io_data_1_out_bits(PE_401_io_data_1_out_bits),
    .io_data_0_in_valid(PE_401_io_data_0_in_valid),
    .io_data_0_in_bits(PE_401_io_data_0_in_bits),
    .io_data_0_out_valid(PE_401_io_data_0_out_valid),
    .io_data_0_out_bits(PE_401_io_data_0_out_bits)
  );
  PE PE_402 ( // @[pe.scala 187:13]
    .clock(PE_402_clock),
    .reset(PE_402_reset),
    .io_data_2_out_valid(PE_402_io_data_2_out_valid),
    .io_data_2_out_bits(PE_402_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_402_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_402_io_data_1_in_valid),
    .io_data_1_in_bits(PE_402_io_data_1_in_bits),
    .io_data_1_out_valid(PE_402_io_data_1_out_valid),
    .io_data_1_out_bits(PE_402_io_data_1_out_bits),
    .io_data_0_in_valid(PE_402_io_data_0_in_valid),
    .io_data_0_in_bits(PE_402_io_data_0_in_bits),
    .io_data_0_out_valid(PE_402_io_data_0_out_valid),
    .io_data_0_out_bits(PE_402_io_data_0_out_bits)
  );
  PE PE_403 ( // @[pe.scala 187:13]
    .clock(PE_403_clock),
    .reset(PE_403_reset),
    .io_data_2_out_valid(PE_403_io_data_2_out_valid),
    .io_data_2_out_bits(PE_403_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_403_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_403_io_data_1_in_valid),
    .io_data_1_in_bits(PE_403_io_data_1_in_bits),
    .io_data_1_out_valid(PE_403_io_data_1_out_valid),
    .io_data_1_out_bits(PE_403_io_data_1_out_bits),
    .io_data_0_in_valid(PE_403_io_data_0_in_valid),
    .io_data_0_in_bits(PE_403_io_data_0_in_bits),
    .io_data_0_out_valid(PE_403_io_data_0_out_valid),
    .io_data_0_out_bits(PE_403_io_data_0_out_bits)
  );
  PE PE_404 ( // @[pe.scala 187:13]
    .clock(PE_404_clock),
    .reset(PE_404_reset),
    .io_data_2_out_valid(PE_404_io_data_2_out_valid),
    .io_data_2_out_bits(PE_404_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_404_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_404_io_data_1_in_valid),
    .io_data_1_in_bits(PE_404_io_data_1_in_bits),
    .io_data_1_out_valid(PE_404_io_data_1_out_valid),
    .io_data_1_out_bits(PE_404_io_data_1_out_bits),
    .io_data_0_in_valid(PE_404_io_data_0_in_valid),
    .io_data_0_in_bits(PE_404_io_data_0_in_bits),
    .io_data_0_out_valid(PE_404_io_data_0_out_valid),
    .io_data_0_out_bits(PE_404_io_data_0_out_bits)
  );
  PE PE_405 ( // @[pe.scala 187:13]
    .clock(PE_405_clock),
    .reset(PE_405_reset),
    .io_data_2_out_valid(PE_405_io_data_2_out_valid),
    .io_data_2_out_bits(PE_405_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_405_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_405_io_data_1_in_valid),
    .io_data_1_in_bits(PE_405_io_data_1_in_bits),
    .io_data_1_out_valid(PE_405_io_data_1_out_valid),
    .io_data_1_out_bits(PE_405_io_data_1_out_bits),
    .io_data_0_in_valid(PE_405_io_data_0_in_valid),
    .io_data_0_in_bits(PE_405_io_data_0_in_bits),
    .io_data_0_out_valid(PE_405_io_data_0_out_valid),
    .io_data_0_out_bits(PE_405_io_data_0_out_bits)
  );
  PE PE_406 ( // @[pe.scala 187:13]
    .clock(PE_406_clock),
    .reset(PE_406_reset),
    .io_data_2_out_valid(PE_406_io_data_2_out_valid),
    .io_data_2_out_bits(PE_406_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_406_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_406_io_data_1_in_valid),
    .io_data_1_in_bits(PE_406_io_data_1_in_bits),
    .io_data_1_out_valid(PE_406_io_data_1_out_valid),
    .io_data_1_out_bits(PE_406_io_data_1_out_bits),
    .io_data_0_in_valid(PE_406_io_data_0_in_valid),
    .io_data_0_in_bits(PE_406_io_data_0_in_bits),
    .io_data_0_out_valid(PE_406_io_data_0_out_valid),
    .io_data_0_out_bits(PE_406_io_data_0_out_bits)
  );
  PE PE_407 ( // @[pe.scala 187:13]
    .clock(PE_407_clock),
    .reset(PE_407_reset),
    .io_data_2_out_valid(PE_407_io_data_2_out_valid),
    .io_data_2_out_bits(PE_407_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_407_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_407_io_data_1_in_valid),
    .io_data_1_in_bits(PE_407_io_data_1_in_bits),
    .io_data_1_out_valid(PE_407_io_data_1_out_valid),
    .io_data_1_out_bits(PE_407_io_data_1_out_bits),
    .io_data_0_in_valid(PE_407_io_data_0_in_valid),
    .io_data_0_in_bits(PE_407_io_data_0_in_bits),
    .io_data_0_out_valid(PE_407_io_data_0_out_valid),
    .io_data_0_out_bits(PE_407_io_data_0_out_bits)
  );
  PE PE_408 ( // @[pe.scala 187:13]
    .clock(PE_408_clock),
    .reset(PE_408_reset),
    .io_data_2_out_valid(PE_408_io_data_2_out_valid),
    .io_data_2_out_bits(PE_408_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_408_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_408_io_data_1_in_valid),
    .io_data_1_in_bits(PE_408_io_data_1_in_bits),
    .io_data_1_out_valid(PE_408_io_data_1_out_valid),
    .io_data_1_out_bits(PE_408_io_data_1_out_bits),
    .io_data_0_in_valid(PE_408_io_data_0_in_valid),
    .io_data_0_in_bits(PE_408_io_data_0_in_bits),
    .io_data_0_out_valid(PE_408_io_data_0_out_valid),
    .io_data_0_out_bits(PE_408_io_data_0_out_bits)
  );
  PE PE_409 ( // @[pe.scala 187:13]
    .clock(PE_409_clock),
    .reset(PE_409_reset),
    .io_data_2_out_valid(PE_409_io_data_2_out_valid),
    .io_data_2_out_bits(PE_409_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_409_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_409_io_data_1_in_valid),
    .io_data_1_in_bits(PE_409_io_data_1_in_bits),
    .io_data_1_out_valid(PE_409_io_data_1_out_valid),
    .io_data_1_out_bits(PE_409_io_data_1_out_bits),
    .io_data_0_in_valid(PE_409_io_data_0_in_valid),
    .io_data_0_in_bits(PE_409_io_data_0_in_bits),
    .io_data_0_out_valid(PE_409_io_data_0_out_valid),
    .io_data_0_out_bits(PE_409_io_data_0_out_bits)
  );
  PE PE_410 ( // @[pe.scala 187:13]
    .clock(PE_410_clock),
    .reset(PE_410_reset),
    .io_data_2_out_valid(PE_410_io_data_2_out_valid),
    .io_data_2_out_bits(PE_410_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_410_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_410_io_data_1_in_valid),
    .io_data_1_in_bits(PE_410_io_data_1_in_bits),
    .io_data_1_out_valid(PE_410_io_data_1_out_valid),
    .io_data_1_out_bits(PE_410_io_data_1_out_bits),
    .io_data_0_in_valid(PE_410_io_data_0_in_valid),
    .io_data_0_in_bits(PE_410_io_data_0_in_bits),
    .io_data_0_out_valid(PE_410_io_data_0_out_valid),
    .io_data_0_out_bits(PE_410_io_data_0_out_bits)
  );
  PE PE_411 ( // @[pe.scala 187:13]
    .clock(PE_411_clock),
    .reset(PE_411_reset),
    .io_data_2_out_valid(PE_411_io_data_2_out_valid),
    .io_data_2_out_bits(PE_411_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_411_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_411_io_data_1_in_valid),
    .io_data_1_in_bits(PE_411_io_data_1_in_bits),
    .io_data_1_out_valid(PE_411_io_data_1_out_valid),
    .io_data_1_out_bits(PE_411_io_data_1_out_bits),
    .io_data_0_in_valid(PE_411_io_data_0_in_valid),
    .io_data_0_in_bits(PE_411_io_data_0_in_bits),
    .io_data_0_out_valid(PE_411_io_data_0_out_valid),
    .io_data_0_out_bits(PE_411_io_data_0_out_bits)
  );
  PE PE_412 ( // @[pe.scala 187:13]
    .clock(PE_412_clock),
    .reset(PE_412_reset),
    .io_data_2_out_valid(PE_412_io_data_2_out_valid),
    .io_data_2_out_bits(PE_412_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_412_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_412_io_data_1_in_valid),
    .io_data_1_in_bits(PE_412_io_data_1_in_bits),
    .io_data_1_out_valid(PE_412_io_data_1_out_valid),
    .io_data_1_out_bits(PE_412_io_data_1_out_bits),
    .io_data_0_in_valid(PE_412_io_data_0_in_valid),
    .io_data_0_in_bits(PE_412_io_data_0_in_bits),
    .io_data_0_out_valid(PE_412_io_data_0_out_valid),
    .io_data_0_out_bits(PE_412_io_data_0_out_bits)
  );
  PE PE_413 ( // @[pe.scala 187:13]
    .clock(PE_413_clock),
    .reset(PE_413_reset),
    .io_data_2_out_valid(PE_413_io_data_2_out_valid),
    .io_data_2_out_bits(PE_413_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_413_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_413_io_data_1_in_valid),
    .io_data_1_in_bits(PE_413_io_data_1_in_bits),
    .io_data_1_out_valid(PE_413_io_data_1_out_valid),
    .io_data_1_out_bits(PE_413_io_data_1_out_bits),
    .io_data_0_in_valid(PE_413_io_data_0_in_valid),
    .io_data_0_in_bits(PE_413_io_data_0_in_bits),
    .io_data_0_out_valid(PE_413_io_data_0_out_valid),
    .io_data_0_out_bits(PE_413_io_data_0_out_bits)
  );
  PE PE_414 ( // @[pe.scala 187:13]
    .clock(PE_414_clock),
    .reset(PE_414_reset),
    .io_data_2_out_valid(PE_414_io_data_2_out_valid),
    .io_data_2_out_bits(PE_414_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_414_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_414_io_data_1_in_valid),
    .io_data_1_in_bits(PE_414_io_data_1_in_bits),
    .io_data_1_out_valid(PE_414_io_data_1_out_valid),
    .io_data_1_out_bits(PE_414_io_data_1_out_bits),
    .io_data_0_in_valid(PE_414_io_data_0_in_valid),
    .io_data_0_in_bits(PE_414_io_data_0_in_bits),
    .io_data_0_out_valid(PE_414_io_data_0_out_valid),
    .io_data_0_out_bits(PE_414_io_data_0_out_bits)
  );
  PE PE_415 ( // @[pe.scala 187:13]
    .clock(PE_415_clock),
    .reset(PE_415_reset),
    .io_data_2_out_valid(PE_415_io_data_2_out_valid),
    .io_data_2_out_bits(PE_415_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_415_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_415_io_data_1_in_valid),
    .io_data_1_in_bits(PE_415_io_data_1_in_bits),
    .io_data_1_out_valid(PE_415_io_data_1_out_valid),
    .io_data_1_out_bits(PE_415_io_data_1_out_bits),
    .io_data_0_in_valid(PE_415_io_data_0_in_valid),
    .io_data_0_in_bits(PE_415_io_data_0_in_bits),
    .io_data_0_out_valid(PE_415_io_data_0_out_valid),
    .io_data_0_out_bits(PE_415_io_data_0_out_bits)
  );
  PE PE_416 ( // @[pe.scala 187:13]
    .clock(PE_416_clock),
    .reset(PE_416_reset),
    .io_data_2_out_valid(PE_416_io_data_2_out_valid),
    .io_data_2_out_bits(PE_416_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_416_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_416_io_data_1_in_valid),
    .io_data_1_in_bits(PE_416_io_data_1_in_bits),
    .io_data_1_out_valid(PE_416_io_data_1_out_valid),
    .io_data_1_out_bits(PE_416_io_data_1_out_bits),
    .io_data_0_in_valid(PE_416_io_data_0_in_valid),
    .io_data_0_in_bits(PE_416_io_data_0_in_bits),
    .io_data_0_out_valid(PE_416_io_data_0_out_valid),
    .io_data_0_out_bits(PE_416_io_data_0_out_bits)
  );
  PE PE_417 ( // @[pe.scala 187:13]
    .clock(PE_417_clock),
    .reset(PE_417_reset),
    .io_data_2_out_valid(PE_417_io_data_2_out_valid),
    .io_data_2_out_bits(PE_417_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_417_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_417_io_data_1_in_valid),
    .io_data_1_in_bits(PE_417_io_data_1_in_bits),
    .io_data_1_out_valid(PE_417_io_data_1_out_valid),
    .io_data_1_out_bits(PE_417_io_data_1_out_bits),
    .io_data_0_in_valid(PE_417_io_data_0_in_valid),
    .io_data_0_in_bits(PE_417_io_data_0_in_bits),
    .io_data_0_out_valid(PE_417_io_data_0_out_valid),
    .io_data_0_out_bits(PE_417_io_data_0_out_bits)
  );
  PE PE_418 ( // @[pe.scala 187:13]
    .clock(PE_418_clock),
    .reset(PE_418_reset),
    .io_data_2_out_valid(PE_418_io_data_2_out_valid),
    .io_data_2_out_bits(PE_418_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_418_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_418_io_data_1_in_valid),
    .io_data_1_in_bits(PE_418_io_data_1_in_bits),
    .io_data_1_out_valid(PE_418_io_data_1_out_valid),
    .io_data_1_out_bits(PE_418_io_data_1_out_bits),
    .io_data_0_in_valid(PE_418_io_data_0_in_valid),
    .io_data_0_in_bits(PE_418_io_data_0_in_bits),
    .io_data_0_out_valid(PE_418_io_data_0_out_valid),
    .io_data_0_out_bits(PE_418_io_data_0_out_bits)
  );
  PE PE_419 ( // @[pe.scala 187:13]
    .clock(PE_419_clock),
    .reset(PE_419_reset),
    .io_data_2_out_valid(PE_419_io_data_2_out_valid),
    .io_data_2_out_bits(PE_419_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_419_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_419_io_data_1_in_valid),
    .io_data_1_in_bits(PE_419_io_data_1_in_bits),
    .io_data_1_out_valid(PE_419_io_data_1_out_valid),
    .io_data_1_out_bits(PE_419_io_data_1_out_bits),
    .io_data_0_in_valid(PE_419_io_data_0_in_valid),
    .io_data_0_in_bits(PE_419_io_data_0_in_bits),
    .io_data_0_out_valid(PE_419_io_data_0_out_valid),
    .io_data_0_out_bits(PE_419_io_data_0_out_bits)
  );
  PE PE_420 ( // @[pe.scala 187:13]
    .clock(PE_420_clock),
    .reset(PE_420_reset),
    .io_data_2_out_valid(PE_420_io_data_2_out_valid),
    .io_data_2_out_bits(PE_420_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_420_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_420_io_data_1_in_valid),
    .io_data_1_in_bits(PE_420_io_data_1_in_bits),
    .io_data_1_out_valid(PE_420_io_data_1_out_valid),
    .io_data_1_out_bits(PE_420_io_data_1_out_bits),
    .io_data_0_in_valid(PE_420_io_data_0_in_valid),
    .io_data_0_in_bits(PE_420_io_data_0_in_bits),
    .io_data_0_out_valid(PE_420_io_data_0_out_valid),
    .io_data_0_out_bits(PE_420_io_data_0_out_bits)
  );
  PE PE_421 ( // @[pe.scala 187:13]
    .clock(PE_421_clock),
    .reset(PE_421_reset),
    .io_data_2_out_valid(PE_421_io_data_2_out_valid),
    .io_data_2_out_bits(PE_421_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_421_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_421_io_data_1_in_valid),
    .io_data_1_in_bits(PE_421_io_data_1_in_bits),
    .io_data_1_out_valid(PE_421_io_data_1_out_valid),
    .io_data_1_out_bits(PE_421_io_data_1_out_bits),
    .io_data_0_in_valid(PE_421_io_data_0_in_valid),
    .io_data_0_in_bits(PE_421_io_data_0_in_bits),
    .io_data_0_out_valid(PE_421_io_data_0_out_valid),
    .io_data_0_out_bits(PE_421_io_data_0_out_bits)
  );
  PE PE_422 ( // @[pe.scala 187:13]
    .clock(PE_422_clock),
    .reset(PE_422_reset),
    .io_data_2_out_valid(PE_422_io_data_2_out_valid),
    .io_data_2_out_bits(PE_422_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_422_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_422_io_data_1_in_valid),
    .io_data_1_in_bits(PE_422_io_data_1_in_bits),
    .io_data_1_out_valid(PE_422_io_data_1_out_valid),
    .io_data_1_out_bits(PE_422_io_data_1_out_bits),
    .io_data_0_in_valid(PE_422_io_data_0_in_valid),
    .io_data_0_in_bits(PE_422_io_data_0_in_bits),
    .io_data_0_out_valid(PE_422_io_data_0_out_valid),
    .io_data_0_out_bits(PE_422_io_data_0_out_bits)
  );
  PE PE_423 ( // @[pe.scala 187:13]
    .clock(PE_423_clock),
    .reset(PE_423_reset),
    .io_data_2_out_valid(PE_423_io_data_2_out_valid),
    .io_data_2_out_bits(PE_423_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_423_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_423_io_data_1_in_valid),
    .io_data_1_in_bits(PE_423_io_data_1_in_bits),
    .io_data_1_out_valid(PE_423_io_data_1_out_valid),
    .io_data_1_out_bits(PE_423_io_data_1_out_bits),
    .io_data_0_in_valid(PE_423_io_data_0_in_valid),
    .io_data_0_in_bits(PE_423_io_data_0_in_bits),
    .io_data_0_out_valid(PE_423_io_data_0_out_valid),
    .io_data_0_out_bits(PE_423_io_data_0_out_bits)
  );
  PE PE_424 ( // @[pe.scala 187:13]
    .clock(PE_424_clock),
    .reset(PE_424_reset),
    .io_data_2_out_valid(PE_424_io_data_2_out_valid),
    .io_data_2_out_bits(PE_424_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_424_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_424_io_data_1_in_valid),
    .io_data_1_in_bits(PE_424_io_data_1_in_bits),
    .io_data_1_out_valid(PE_424_io_data_1_out_valid),
    .io_data_1_out_bits(PE_424_io_data_1_out_bits),
    .io_data_0_in_valid(PE_424_io_data_0_in_valid),
    .io_data_0_in_bits(PE_424_io_data_0_in_bits),
    .io_data_0_out_valid(PE_424_io_data_0_out_valid),
    .io_data_0_out_bits(PE_424_io_data_0_out_bits)
  );
  PE PE_425 ( // @[pe.scala 187:13]
    .clock(PE_425_clock),
    .reset(PE_425_reset),
    .io_data_2_out_valid(PE_425_io_data_2_out_valid),
    .io_data_2_out_bits(PE_425_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_425_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_425_io_data_1_in_valid),
    .io_data_1_in_bits(PE_425_io_data_1_in_bits),
    .io_data_1_out_valid(PE_425_io_data_1_out_valid),
    .io_data_1_out_bits(PE_425_io_data_1_out_bits),
    .io_data_0_in_valid(PE_425_io_data_0_in_valid),
    .io_data_0_in_bits(PE_425_io_data_0_in_bits),
    .io_data_0_out_valid(PE_425_io_data_0_out_valid),
    .io_data_0_out_bits(PE_425_io_data_0_out_bits)
  );
  PE PE_426 ( // @[pe.scala 187:13]
    .clock(PE_426_clock),
    .reset(PE_426_reset),
    .io_data_2_out_valid(PE_426_io_data_2_out_valid),
    .io_data_2_out_bits(PE_426_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_426_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_426_io_data_1_in_valid),
    .io_data_1_in_bits(PE_426_io_data_1_in_bits),
    .io_data_1_out_valid(PE_426_io_data_1_out_valid),
    .io_data_1_out_bits(PE_426_io_data_1_out_bits),
    .io_data_0_in_valid(PE_426_io_data_0_in_valid),
    .io_data_0_in_bits(PE_426_io_data_0_in_bits),
    .io_data_0_out_valid(PE_426_io_data_0_out_valid),
    .io_data_0_out_bits(PE_426_io_data_0_out_bits)
  );
  PE PE_427 ( // @[pe.scala 187:13]
    .clock(PE_427_clock),
    .reset(PE_427_reset),
    .io_data_2_out_valid(PE_427_io_data_2_out_valid),
    .io_data_2_out_bits(PE_427_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_427_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_427_io_data_1_in_valid),
    .io_data_1_in_bits(PE_427_io_data_1_in_bits),
    .io_data_1_out_valid(PE_427_io_data_1_out_valid),
    .io_data_1_out_bits(PE_427_io_data_1_out_bits),
    .io_data_0_in_valid(PE_427_io_data_0_in_valid),
    .io_data_0_in_bits(PE_427_io_data_0_in_bits),
    .io_data_0_out_valid(PE_427_io_data_0_out_valid),
    .io_data_0_out_bits(PE_427_io_data_0_out_bits)
  );
  PE PE_428 ( // @[pe.scala 187:13]
    .clock(PE_428_clock),
    .reset(PE_428_reset),
    .io_data_2_out_valid(PE_428_io_data_2_out_valid),
    .io_data_2_out_bits(PE_428_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_428_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_428_io_data_1_in_valid),
    .io_data_1_in_bits(PE_428_io_data_1_in_bits),
    .io_data_1_out_valid(PE_428_io_data_1_out_valid),
    .io_data_1_out_bits(PE_428_io_data_1_out_bits),
    .io_data_0_in_valid(PE_428_io_data_0_in_valid),
    .io_data_0_in_bits(PE_428_io_data_0_in_bits),
    .io_data_0_out_valid(PE_428_io_data_0_out_valid),
    .io_data_0_out_bits(PE_428_io_data_0_out_bits)
  );
  PE PE_429 ( // @[pe.scala 187:13]
    .clock(PE_429_clock),
    .reset(PE_429_reset),
    .io_data_2_out_valid(PE_429_io_data_2_out_valid),
    .io_data_2_out_bits(PE_429_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_429_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_429_io_data_1_in_valid),
    .io_data_1_in_bits(PE_429_io_data_1_in_bits),
    .io_data_1_out_valid(PE_429_io_data_1_out_valid),
    .io_data_1_out_bits(PE_429_io_data_1_out_bits),
    .io_data_0_in_valid(PE_429_io_data_0_in_valid),
    .io_data_0_in_bits(PE_429_io_data_0_in_bits),
    .io_data_0_out_valid(PE_429_io_data_0_out_valid),
    .io_data_0_out_bits(PE_429_io_data_0_out_bits)
  );
  PE PE_430 ( // @[pe.scala 187:13]
    .clock(PE_430_clock),
    .reset(PE_430_reset),
    .io_data_2_out_valid(PE_430_io_data_2_out_valid),
    .io_data_2_out_bits(PE_430_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_430_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_430_io_data_1_in_valid),
    .io_data_1_in_bits(PE_430_io_data_1_in_bits),
    .io_data_1_out_valid(PE_430_io_data_1_out_valid),
    .io_data_1_out_bits(PE_430_io_data_1_out_bits),
    .io_data_0_in_valid(PE_430_io_data_0_in_valid),
    .io_data_0_in_bits(PE_430_io_data_0_in_bits),
    .io_data_0_out_valid(PE_430_io_data_0_out_valid),
    .io_data_0_out_bits(PE_430_io_data_0_out_bits)
  );
  PE PE_431 ( // @[pe.scala 187:13]
    .clock(PE_431_clock),
    .reset(PE_431_reset),
    .io_data_2_out_valid(PE_431_io_data_2_out_valid),
    .io_data_2_out_bits(PE_431_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_431_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_431_io_data_1_in_valid),
    .io_data_1_in_bits(PE_431_io_data_1_in_bits),
    .io_data_1_out_valid(PE_431_io_data_1_out_valid),
    .io_data_1_out_bits(PE_431_io_data_1_out_bits),
    .io_data_0_in_valid(PE_431_io_data_0_in_valid),
    .io_data_0_in_bits(PE_431_io_data_0_in_bits),
    .io_data_0_out_valid(PE_431_io_data_0_out_valid),
    .io_data_0_out_bits(PE_431_io_data_0_out_bits)
  );
  PE PE_432 ( // @[pe.scala 187:13]
    .clock(PE_432_clock),
    .reset(PE_432_reset),
    .io_data_2_out_valid(PE_432_io_data_2_out_valid),
    .io_data_2_out_bits(PE_432_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_432_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_432_io_data_1_in_valid),
    .io_data_1_in_bits(PE_432_io_data_1_in_bits),
    .io_data_1_out_valid(PE_432_io_data_1_out_valid),
    .io_data_1_out_bits(PE_432_io_data_1_out_bits),
    .io_data_0_in_valid(PE_432_io_data_0_in_valid),
    .io_data_0_in_bits(PE_432_io_data_0_in_bits),
    .io_data_0_out_valid(PE_432_io_data_0_out_valid),
    .io_data_0_out_bits(PE_432_io_data_0_out_bits)
  );
  PE PE_433 ( // @[pe.scala 187:13]
    .clock(PE_433_clock),
    .reset(PE_433_reset),
    .io_data_2_out_valid(PE_433_io_data_2_out_valid),
    .io_data_2_out_bits(PE_433_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_433_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_433_io_data_1_in_valid),
    .io_data_1_in_bits(PE_433_io_data_1_in_bits),
    .io_data_1_out_valid(PE_433_io_data_1_out_valid),
    .io_data_1_out_bits(PE_433_io_data_1_out_bits),
    .io_data_0_in_valid(PE_433_io_data_0_in_valid),
    .io_data_0_in_bits(PE_433_io_data_0_in_bits),
    .io_data_0_out_valid(PE_433_io_data_0_out_valid),
    .io_data_0_out_bits(PE_433_io_data_0_out_bits)
  );
  PE PE_434 ( // @[pe.scala 187:13]
    .clock(PE_434_clock),
    .reset(PE_434_reset),
    .io_data_2_out_valid(PE_434_io_data_2_out_valid),
    .io_data_2_out_bits(PE_434_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_434_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_434_io_data_1_in_valid),
    .io_data_1_in_bits(PE_434_io_data_1_in_bits),
    .io_data_1_out_valid(PE_434_io_data_1_out_valid),
    .io_data_1_out_bits(PE_434_io_data_1_out_bits),
    .io_data_0_in_valid(PE_434_io_data_0_in_valid),
    .io_data_0_in_bits(PE_434_io_data_0_in_bits),
    .io_data_0_out_valid(PE_434_io_data_0_out_valid),
    .io_data_0_out_bits(PE_434_io_data_0_out_bits)
  );
  PE PE_435 ( // @[pe.scala 187:13]
    .clock(PE_435_clock),
    .reset(PE_435_reset),
    .io_data_2_out_valid(PE_435_io_data_2_out_valid),
    .io_data_2_out_bits(PE_435_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_435_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_435_io_data_1_in_valid),
    .io_data_1_in_bits(PE_435_io_data_1_in_bits),
    .io_data_1_out_valid(PE_435_io_data_1_out_valid),
    .io_data_1_out_bits(PE_435_io_data_1_out_bits),
    .io_data_0_in_valid(PE_435_io_data_0_in_valid),
    .io_data_0_in_bits(PE_435_io_data_0_in_bits),
    .io_data_0_out_valid(PE_435_io_data_0_out_valid),
    .io_data_0_out_bits(PE_435_io_data_0_out_bits)
  );
  PE PE_436 ( // @[pe.scala 187:13]
    .clock(PE_436_clock),
    .reset(PE_436_reset),
    .io_data_2_out_valid(PE_436_io_data_2_out_valid),
    .io_data_2_out_bits(PE_436_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_436_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_436_io_data_1_in_valid),
    .io_data_1_in_bits(PE_436_io_data_1_in_bits),
    .io_data_1_out_valid(PE_436_io_data_1_out_valid),
    .io_data_1_out_bits(PE_436_io_data_1_out_bits),
    .io_data_0_in_valid(PE_436_io_data_0_in_valid),
    .io_data_0_in_bits(PE_436_io_data_0_in_bits),
    .io_data_0_out_valid(PE_436_io_data_0_out_valid),
    .io_data_0_out_bits(PE_436_io_data_0_out_bits)
  );
  PE PE_437 ( // @[pe.scala 187:13]
    .clock(PE_437_clock),
    .reset(PE_437_reset),
    .io_data_2_out_valid(PE_437_io_data_2_out_valid),
    .io_data_2_out_bits(PE_437_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_437_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_437_io_data_1_in_valid),
    .io_data_1_in_bits(PE_437_io_data_1_in_bits),
    .io_data_1_out_valid(PE_437_io_data_1_out_valid),
    .io_data_1_out_bits(PE_437_io_data_1_out_bits),
    .io_data_0_in_valid(PE_437_io_data_0_in_valid),
    .io_data_0_in_bits(PE_437_io_data_0_in_bits),
    .io_data_0_out_valid(PE_437_io_data_0_out_valid),
    .io_data_0_out_bits(PE_437_io_data_0_out_bits)
  );
  PE PE_438 ( // @[pe.scala 187:13]
    .clock(PE_438_clock),
    .reset(PE_438_reset),
    .io_data_2_out_valid(PE_438_io_data_2_out_valid),
    .io_data_2_out_bits(PE_438_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_438_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_438_io_data_1_in_valid),
    .io_data_1_in_bits(PE_438_io_data_1_in_bits),
    .io_data_1_out_valid(PE_438_io_data_1_out_valid),
    .io_data_1_out_bits(PE_438_io_data_1_out_bits),
    .io_data_0_in_valid(PE_438_io_data_0_in_valid),
    .io_data_0_in_bits(PE_438_io_data_0_in_bits),
    .io_data_0_out_valid(PE_438_io_data_0_out_valid),
    .io_data_0_out_bits(PE_438_io_data_0_out_bits)
  );
  PE PE_439 ( // @[pe.scala 187:13]
    .clock(PE_439_clock),
    .reset(PE_439_reset),
    .io_data_2_out_valid(PE_439_io_data_2_out_valid),
    .io_data_2_out_bits(PE_439_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_439_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_439_io_data_1_in_valid),
    .io_data_1_in_bits(PE_439_io_data_1_in_bits),
    .io_data_1_out_valid(PE_439_io_data_1_out_valid),
    .io_data_1_out_bits(PE_439_io_data_1_out_bits),
    .io_data_0_in_valid(PE_439_io_data_0_in_valid),
    .io_data_0_in_bits(PE_439_io_data_0_in_bits),
    .io_data_0_out_valid(PE_439_io_data_0_out_valid),
    .io_data_0_out_bits(PE_439_io_data_0_out_bits)
  );
  PE PE_440 ( // @[pe.scala 187:13]
    .clock(PE_440_clock),
    .reset(PE_440_reset),
    .io_data_2_out_valid(PE_440_io_data_2_out_valid),
    .io_data_2_out_bits(PE_440_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_440_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_440_io_data_1_in_valid),
    .io_data_1_in_bits(PE_440_io_data_1_in_bits),
    .io_data_1_out_valid(PE_440_io_data_1_out_valid),
    .io_data_1_out_bits(PE_440_io_data_1_out_bits),
    .io_data_0_in_valid(PE_440_io_data_0_in_valid),
    .io_data_0_in_bits(PE_440_io_data_0_in_bits),
    .io_data_0_out_valid(PE_440_io_data_0_out_valid),
    .io_data_0_out_bits(PE_440_io_data_0_out_bits)
  );
  PE PE_441 ( // @[pe.scala 187:13]
    .clock(PE_441_clock),
    .reset(PE_441_reset),
    .io_data_2_out_valid(PE_441_io_data_2_out_valid),
    .io_data_2_out_bits(PE_441_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_441_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_441_io_data_1_in_valid),
    .io_data_1_in_bits(PE_441_io_data_1_in_bits),
    .io_data_1_out_valid(PE_441_io_data_1_out_valid),
    .io_data_1_out_bits(PE_441_io_data_1_out_bits),
    .io_data_0_in_valid(PE_441_io_data_0_in_valid),
    .io_data_0_in_bits(PE_441_io_data_0_in_bits),
    .io_data_0_out_valid(PE_441_io_data_0_out_valid),
    .io_data_0_out_bits(PE_441_io_data_0_out_bits)
  );
  PE PE_442 ( // @[pe.scala 187:13]
    .clock(PE_442_clock),
    .reset(PE_442_reset),
    .io_data_2_out_valid(PE_442_io_data_2_out_valid),
    .io_data_2_out_bits(PE_442_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_442_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_442_io_data_1_in_valid),
    .io_data_1_in_bits(PE_442_io_data_1_in_bits),
    .io_data_1_out_valid(PE_442_io_data_1_out_valid),
    .io_data_1_out_bits(PE_442_io_data_1_out_bits),
    .io_data_0_in_valid(PE_442_io_data_0_in_valid),
    .io_data_0_in_bits(PE_442_io_data_0_in_bits),
    .io_data_0_out_valid(PE_442_io_data_0_out_valid),
    .io_data_0_out_bits(PE_442_io_data_0_out_bits)
  );
  PE PE_443 ( // @[pe.scala 187:13]
    .clock(PE_443_clock),
    .reset(PE_443_reset),
    .io_data_2_out_valid(PE_443_io_data_2_out_valid),
    .io_data_2_out_bits(PE_443_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_443_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_443_io_data_1_in_valid),
    .io_data_1_in_bits(PE_443_io_data_1_in_bits),
    .io_data_1_out_valid(PE_443_io_data_1_out_valid),
    .io_data_1_out_bits(PE_443_io_data_1_out_bits),
    .io_data_0_in_valid(PE_443_io_data_0_in_valid),
    .io_data_0_in_bits(PE_443_io_data_0_in_bits),
    .io_data_0_out_valid(PE_443_io_data_0_out_valid),
    .io_data_0_out_bits(PE_443_io_data_0_out_bits)
  );
  PE PE_444 ( // @[pe.scala 187:13]
    .clock(PE_444_clock),
    .reset(PE_444_reset),
    .io_data_2_out_valid(PE_444_io_data_2_out_valid),
    .io_data_2_out_bits(PE_444_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_444_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_444_io_data_1_in_valid),
    .io_data_1_in_bits(PE_444_io_data_1_in_bits),
    .io_data_1_out_valid(PE_444_io_data_1_out_valid),
    .io_data_1_out_bits(PE_444_io_data_1_out_bits),
    .io_data_0_in_valid(PE_444_io_data_0_in_valid),
    .io_data_0_in_bits(PE_444_io_data_0_in_bits),
    .io_data_0_out_valid(PE_444_io_data_0_out_valid),
    .io_data_0_out_bits(PE_444_io_data_0_out_bits)
  );
  PE PE_445 ( // @[pe.scala 187:13]
    .clock(PE_445_clock),
    .reset(PE_445_reset),
    .io_data_2_out_valid(PE_445_io_data_2_out_valid),
    .io_data_2_out_bits(PE_445_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_445_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_445_io_data_1_in_valid),
    .io_data_1_in_bits(PE_445_io_data_1_in_bits),
    .io_data_1_out_valid(PE_445_io_data_1_out_valid),
    .io_data_1_out_bits(PE_445_io_data_1_out_bits),
    .io_data_0_in_valid(PE_445_io_data_0_in_valid),
    .io_data_0_in_bits(PE_445_io_data_0_in_bits),
    .io_data_0_out_valid(PE_445_io_data_0_out_valid),
    .io_data_0_out_bits(PE_445_io_data_0_out_bits)
  );
  PE PE_446 ( // @[pe.scala 187:13]
    .clock(PE_446_clock),
    .reset(PE_446_reset),
    .io_data_2_out_valid(PE_446_io_data_2_out_valid),
    .io_data_2_out_bits(PE_446_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_446_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_446_io_data_1_in_valid),
    .io_data_1_in_bits(PE_446_io_data_1_in_bits),
    .io_data_1_out_valid(PE_446_io_data_1_out_valid),
    .io_data_1_out_bits(PE_446_io_data_1_out_bits),
    .io_data_0_in_valid(PE_446_io_data_0_in_valid),
    .io_data_0_in_bits(PE_446_io_data_0_in_bits),
    .io_data_0_out_valid(PE_446_io_data_0_out_valid),
    .io_data_0_out_bits(PE_446_io_data_0_out_bits)
  );
  PE PE_447 ( // @[pe.scala 187:13]
    .clock(PE_447_clock),
    .reset(PE_447_reset),
    .io_data_2_out_valid(PE_447_io_data_2_out_valid),
    .io_data_2_out_bits(PE_447_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_447_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_447_io_data_1_in_valid),
    .io_data_1_in_bits(PE_447_io_data_1_in_bits),
    .io_data_1_out_valid(PE_447_io_data_1_out_valid),
    .io_data_1_out_bits(PE_447_io_data_1_out_bits),
    .io_data_0_in_valid(PE_447_io_data_0_in_valid),
    .io_data_0_in_bits(PE_447_io_data_0_in_bits),
    .io_data_0_out_valid(PE_447_io_data_0_out_valid),
    .io_data_0_out_bits(PE_447_io_data_0_out_bits)
  );
  PE PE_448 ( // @[pe.scala 187:13]
    .clock(PE_448_clock),
    .reset(PE_448_reset),
    .io_data_2_out_valid(PE_448_io_data_2_out_valid),
    .io_data_2_out_bits(PE_448_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_448_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_448_io_data_1_in_valid),
    .io_data_1_in_bits(PE_448_io_data_1_in_bits),
    .io_data_1_out_valid(PE_448_io_data_1_out_valid),
    .io_data_1_out_bits(PE_448_io_data_1_out_bits),
    .io_data_0_in_valid(PE_448_io_data_0_in_valid),
    .io_data_0_in_bits(PE_448_io_data_0_in_bits),
    .io_data_0_out_valid(PE_448_io_data_0_out_valid),
    .io_data_0_out_bits(PE_448_io_data_0_out_bits)
  );
  PE PE_449 ( // @[pe.scala 187:13]
    .clock(PE_449_clock),
    .reset(PE_449_reset),
    .io_data_2_out_valid(PE_449_io_data_2_out_valid),
    .io_data_2_out_bits(PE_449_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_449_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_449_io_data_1_in_valid),
    .io_data_1_in_bits(PE_449_io_data_1_in_bits),
    .io_data_1_out_valid(PE_449_io_data_1_out_valid),
    .io_data_1_out_bits(PE_449_io_data_1_out_bits),
    .io_data_0_in_valid(PE_449_io_data_0_in_valid),
    .io_data_0_in_bits(PE_449_io_data_0_in_bits),
    .io_data_0_out_valid(PE_449_io_data_0_out_valid),
    .io_data_0_out_bits(PE_449_io_data_0_out_bits)
  );
  PE PE_450 ( // @[pe.scala 187:13]
    .clock(PE_450_clock),
    .reset(PE_450_reset),
    .io_data_2_out_valid(PE_450_io_data_2_out_valid),
    .io_data_2_out_bits(PE_450_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_450_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_450_io_data_1_in_valid),
    .io_data_1_in_bits(PE_450_io_data_1_in_bits),
    .io_data_1_out_valid(PE_450_io_data_1_out_valid),
    .io_data_1_out_bits(PE_450_io_data_1_out_bits),
    .io_data_0_in_valid(PE_450_io_data_0_in_valid),
    .io_data_0_in_bits(PE_450_io_data_0_in_bits),
    .io_data_0_out_valid(PE_450_io_data_0_out_valid),
    .io_data_0_out_bits(PE_450_io_data_0_out_bits)
  );
  PE PE_451 ( // @[pe.scala 187:13]
    .clock(PE_451_clock),
    .reset(PE_451_reset),
    .io_data_2_out_valid(PE_451_io_data_2_out_valid),
    .io_data_2_out_bits(PE_451_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_451_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_451_io_data_1_in_valid),
    .io_data_1_in_bits(PE_451_io_data_1_in_bits),
    .io_data_1_out_valid(PE_451_io_data_1_out_valid),
    .io_data_1_out_bits(PE_451_io_data_1_out_bits),
    .io_data_0_in_valid(PE_451_io_data_0_in_valid),
    .io_data_0_in_bits(PE_451_io_data_0_in_bits),
    .io_data_0_out_valid(PE_451_io_data_0_out_valid),
    .io_data_0_out_bits(PE_451_io_data_0_out_bits)
  );
  PE PE_452 ( // @[pe.scala 187:13]
    .clock(PE_452_clock),
    .reset(PE_452_reset),
    .io_data_2_out_valid(PE_452_io_data_2_out_valid),
    .io_data_2_out_bits(PE_452_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_452_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_452_io_data_1_in_valid),
    .io_data_1_in_bits(PE_452_io_data_1_in_bits),
    .io_data_1_out_valid(PE_452_io_data_1_out_valid),
    .io_data_1_out_bits(PE_452_io_data_1_out_bits),
    .io_data_0_in_valid(PE_452_io_data_0_in_valid),
    .io_data_0_in_bits(PE_452_io_data_0_in_bits),
    .io_data_0_out_valid(PE_452_io_data_0_out_valid),
    .io_data_0_out_bits(PE_452_io_data_0_out_bits)
  );
  PE PE_453 ( // @[pe.scala 187:13]
    .clock(PE_453_clock),
    .reset(PE_453_reset),
    .io_data_2_out_valid(PE_453_io_data_2_out_valid),
    .io_data_2_out_bits(PE_453_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_453_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_453_io_data_1_in_valid),
    .io_data_1_in_bits(PE_453_io_data_1_in_bits),
    .io_data_1_out_valid(PE_453_io_data_1_out_valid),
    .io_data_1_out_bits(PE_453_io_data_1_out_bits),
    .io_data_0_in_valid(PE_453_io_data_0_in_valid),
    .io_data_0_in_bits(PE_453_io_data_0_in_bits),
    .io_data_0_out_valid(PE_453_io_data_0_out_valid),
    .io_data_0_out_bits(PE_453_io_data_0_out_bits)
  );
  PE PE_454 ( // @[pe.scala 187:13]
    .clock(PE_454_clock),
    .reset(PE_454_reset),
    .io_data_2_out_valid(PE_454_io_data_2_out_valid),
    .io_data_2_out_bits(PE_454_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_454_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_454_io_data_1_in_valid),
    .io_data_1_in_bits(PE_454_io_data_1_in_bits),
    .io_data_1_out_valid(PE_454_io_data_1_out_valid),
    .io_data_1_out_bits(PE_454_io_data_1_out_bits),
    .io_data_0_in_valid(PE_454_io_data_0_in_valid),
    .io_data_0_in_bits(PE_454_io_data_0_in_bits),
    .io_data_0_out_valid(PE_454_io_data_0_out_valid),
    .io_data_0_out_bits(PE_454_io_data_0_out_bits)
  );
  PE PE_455 ( // @[pe.scala 187:13]
    .clock(PE_455_clock),
    .reset(PE_455_reset),
    .io_data_2_out_valid(PE_455_io_data_2_out_valid),
    .io_data_2_out_bits(PE_455_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_455_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_455_io_data_1_in_valid),
    .io_data_1_in_bits(PE_455_io_data_1_in_bits),
    .io_data_1_out_valid(PE_455_io_data_1_out_valid),
    .io_data_1_out_bits(PE_455_io_data_1_out_bits),
    .io_data_0_in_valid(PE_455_io_data_0_in_valid),
    .io_data_0_in_bits(PE_455_io_data_0_in_bits),
    .io_data_0_out_valid(PE_455_io_data_0_out_valid),
    .io_data_0_out_bits(PE_455_io_data_0_out_bits)
  );
  PE PE_456 ( // @[pe.scala 187:13]
    .clock(PE_456_clock),
    .reset(PE_456_reset),
    .io_data_2_out_valid(PE_456_io_data_2_out_valid),
    .io_data_2_out_bits(PE_456_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_456_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_456_io_data_1_in_valid),
    .io_data_1_in_bits(PE_456_io_data_1_in_bits),
    .io_data_1_out_valid(PE_456_io_data_1_out_valid),
    .io_data_1_out_bits(PE_456_io_data_1_out_bits),
    .io_data_0_in_valid(PE_456_io_data_0_in_valid),
    .io_data_0_in_bits(PE_456_io_data_0_in_bits),
    .io_data_0_out_valid(PE_456_io_data_0_out_valid),
    .io_data_0_out_bits(PE_456_io_data_0_out_bits)
  );
  PE PE_457 ( // @[pe.scala 187:13]
    .clock(PE_457_clock),
    .reset(PE_457_reset),
    .io_data_2_out_valid(PE_457_io_data_2_out_valid),
    .io_data_2_out_bits(PE_457_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_457_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_457_io_data_1_in_valid),
    .io_data_1_in_bits(PE_457_io_data_1_in_bits),
    .io_data_1_out_valid(PE_457_io_data_1_out_valid),
    .io_data_1_out_bits(PE_457_io_data_1_out_bits),
    .io_data_0_in_valid(PE_457_io_data_0_in_valid),
    .io_data_0_in_bits(PE_457_io_data_0_in_bits),
    .io_data_0_out_valid(PE_457_io_data_0_out_valid),
    .io_data_0_out_bits(PE_457_io_data_0_out_bits)
  );
  PE PE_458 ( // @[pe.scala 187:13]
    .clock(PE_458_clock),
    .reset(PE_458_reset),
    .io_data_2_out_valid(PE_458_io_data_2_out_valid),
    .io_data_2_out_bits(PE_458_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_458_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_458_io_data_1_in_valid),
    .io_data_1_in_bits(PE_458_io_data_1_in_bits),
    .io_data_1_out_valid(PE_458_io_data_1_out_valid),
    .io_data_1_out_bits(PE_458_io_data_1_out_bits),
    .io_data_0_in_valid(PE_458_io_data_0_in_valid),
    .io_data_0_in_bits(PE_458_io_data_0_in_bits),
    .io_data_0_out_valid(PE_458_io_data_0_out_valid),
    .io_data_0_out_bits(PE_458_io_data_0_out_bits)
  );
  PE PE_459 ( // @[pe.scala 187:13]
    .clock(PE_459_clock),
    .reset(PE_459_reset),
    .io_data_2_out_valid(PE_459_io_data_2_out_valid),
    .io_data_2_out_bits(PE_459_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_459_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_459_io_data_1_in_valid),
    .io_data_1_in_bits(PE_459_io_data_1_in_bits),
    .io_data_1_out_valid(PE_459_io_data_1_out_valid),
    .io_data_1_out_bits(PE_459_io_data_1_out_bits),
    .io_data_0_in_valid(PE_459_io_data_0_in_valid),
    .io_data_0_in_bits(PE_459_io_data_0_in_bits),
    .io_data_0_out_valid(PE_459_io_data_0_out_valid),
    .io_data_0_out_bits(PE_459_io_data_0_out_bits)
  );
  PE PE_460 ( // @[pe.scala 187:13]
    .clock(PE_460_clock),
    .reset(PE_460_reset),
    .io_data_2_out_valid(PE_460_io_data_2_out_valid),
    .io_data_2_out_bits(PE_460_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_460_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_460_io_data_1_in_valid),
    .io_data_1_in_bits(PE_460_io_data_1_in_bits),
    .io_data_1_out_valid(PE_460_io_data_1_out_valid),
    .io_data_1_out_bits(PE_460_io_data_1_out_bits),
    .io_data_0_in_valid(PE_460_io_data_0_in_valid),
    .io_data_0_in_bits(PE_460_io_data_0_in_bits),
    .io_data_0_out_valid(PE_460_io_data_0_out_valid),
    .io_data_0_out_bits(PE_460_io_data_0_out_bits)
  );
  PE PE_461 ( // @[pe.scala 187:13]
    .clock(PE_461_clock),
    .reset(PE_461_reset),
    .io_data_2_out_valid(PE_461_io_data_2_out_valid),
    .io_data_2_out_bits(PE_461_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_461_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_461_io_data_1_in_valid),
    .io_data_1_in_bits(PE_461_io_data_1_in_bits),
    .io_data_1_out_valid(PE_461_io_data_1_out_valid),
    .io_data_1_out_bits(PE_461_io_data_1_out_bits),
    .io_data_0_in_valid(PE_461_io_data_0_in_valid),
    .io_data_0_in_bits(PE_461_io_data_0_in_bits),
    .io_data_0_out_valid(PE_461_io_data_0_out_valid),
    .io_data_0_out_bits(PE_461_io_data_0_out_bits)
  );
  PE PE_462 ( // @[pe.scala 187:13]
    .clock(PE_462_clock),
    .reset(PE_462_reset),
    .io_data_2_out_valid(PE_462_io_data_2_out_valid),
    .io_data_2_out_bits(PE_462_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_462_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_462_io_data_1_in_valid),
    .io_data_1_in_bits(PE_462_io_data_1_in_bits),
    .io_data_1_out_valid(PE_462_io_data_1_out_valid),
    .io_data_1_out_bits(PE_462_io_data_1_out_bits),
    .io_data_0_in_valid(PE_462_io_data_0_in_valid),
    .io_data_0_in_bits(PE_462_io_data_0_in_bits),
    .io_data_0_out_valid(PE_462_io_data_0_out_valid),
    .io_data_0_out_bits(PE_462_io_data_0_out_bits)
  );
  PE PE_463 ( // @[pe.scala 187:13]
    .clock(PE_463_clock),
    .reset(PE_463_reset),
    .io_data_2_out_valid(PE_463_io_data_2_out_valid),
    .io_data_2_out_bits(PE_463_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_463_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_463_io_data_1_in_valid),
    .io_data_1_in_bits(PE_463_io_data_1_in_bits),
    .io_data_1_out_valid(PE_463_io_data_1_out_valid),
    .io_data_1_out_bits(PE_463_io_data_1_out_bits),
    .io_data_0_in_valid(PE_463_io_data_0_in_valid),
    .io_data_0_in_bits(PE_463_io_data_0_in_bits),
    .io_data_0_out_valid(PE_463_io_data_0_out_valid),
    .io_data_0_out_bits(PE_463_io_data_0_out_bits)
  );
  PE PE_464 ( // @[pe.scala 187:13]
    .clock(PE_464_clock),
    .reset(PE_464_reset),
    .io_data_2_out_valid(PE_464_io_data_2_out_valid),
    .io_data_2_out_bits(PE_464_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_464_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_464_io_data_1_in_valid),
    .io_data_1_in_bits(PE_464_io_data_1_in_bits),
    .io_data_1_out_valid(PE_464_io_data_1_out_valid),
    .io_data_1_out_bits(PE_464_io_data_1_out_bits),
    .io_data_0_in_valid(PE_464_io_data_0_in_valid),
    .io_data_0_in_bits(PE_464_io_data_0_in_bits),
    .io_data_0_out_valid(PE_464_io_data_0_out_valid),
    .io_data_0_out_bits(PE_464_io_data_0_out_bits)
  );
  PE PE_465 ( // @[pe.scala 187:13]
    .clock(PE_465_clock),
    .reset(PE_465_reset),
    .io_data_2_out_valid(PE_465_io_data_2_out_valid),
    .io_data_2_out_bits(PE_465_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_465_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_465_io_data_1_in_valid),
    .io_data_1_in_bits(PE_465_io_data_1_in_bits),
    .io_data_1_out_valid(PE_465_io_data_1_out_valid),
    .io_data_1_out_bits(PE_465_io_data_1_out_bits),
    .io_data_0_in_valid(PE_465_io_data_0_in_valid),
    .io_data_0_in_bits(PE_465_io_data_0_in_bits),
    .io_data_0_out_valid(PE_465_io_data_0_out_valid),
    .io_data_0_out_bits(PE_465_io_data_0_out_bits)
  );
  PE PE_466 ( // @[pe.scala 187:13]
    .clock(PE_466_clock),
    .reset(PE_466_reset),
    .io_data_2_out_valid(PE_466_io_data_2_out_valid),
    .io_data_2_out_bits(PE_466_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_466_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_466_io_data_1_in_valid),
    .io_data_1_in_bits(PE_466_io_data_1_in_bits),
    .io_data_1_out_valid(PE_466_io_data_1_out_valid),
    .io_data_1_out_bits(PE_466_io_data_1_out_bits),
    .io_data_0_in_valid(PE_466_io_data_0_in_valid),
    .io_data_0_in_bits(PE_466_io_data_0_in_bits),
    .io_data_0_out_valid(PE_466_io_data_0_out_valid),
    .io_data_0_out_bits(PE_466_io_data_0_out_bits)
  );
  PE PE_467 ( // @[pe.scala 187:13]
    .clock(PE_467_clock),
    .reset(PE_467_reset),
    .io_data_2_out_valid(PE_467_io_data_2_out_valid),
    .io_data_2_out_bits(PE_467_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_467_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_467_io_data_1_in_valid),
    .io_data_1_in_bits(PE_467_io_data_1_in_bits),
    .io_data_1_out_valid(PE_467_io_data_1_out_valid),
    .io_data_1_out_bits(PE_467_io_data_1_out_bits),
    .io_data_0_in_valid(PE_467_io_data_0_in_valid),
    .io_data_0_in_bits(PE_467_io_data_0_in_bits),
    .io_data_0_out_valid(PE_467_io_data_0_out_valid),
    .io_data_0_out_bits(PE_467_io_data_0_out_bits)
  );
  PE PE_468 ( // @[pe.scala 187:13]
    .clock(PE_468_clock),
    .reset(PE_468_reset),
    .io_data_2_out_valid(PE_468_io_data_2_out_valid),
    .io_data_2_out_bits(PE_468_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_468_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_468_io_data_1_in_valid),
    .io_data_1_in_bits(PE_468_io_data_1_in_bits),
    .io_data_1_out_valid(PE_468_io_data_1_out_valid),
    .io_data_1_out_bits(PE_468_io_data_1_out_bits),
    .io_data_0_in_valid(PE_468_io_data_0_in_valid),
    .io_data_0_in_bits(PE_468_io_data_0_in_bits),
    .io_data_0_out_valid(PE_468_io_data_0_out_valid),
    .io_data_0_out_bits(PE_468_io_data_0_out_bits)
  );
  PE PE_469 ( // @[pe.scala 187:13]
    .clock(PE_469_clock),
    .reset(PE_469_reset),
    .io_data_2_out_valid(PE_469_io_data_2_out_valid),
    .io_data_2_out_bits(PE_469_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_469_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_469_io_data_1_in_valid),
    .io_data_1_in_bits(PE_469_io_data_1_in_bits),
    .io_data_1_out_valid(PE_469_io_data_1_out_valid),
    .io_data_1_out_bits(PE_469_io_data_1_out_bits),
    .io_data_0_in_valid(PE_469_io_data_0_in_valid),
    .io_data_0_in_bits(PE_469_io_data_0_in_bits),
    .io_data_0_out_valid(PE_469_io_data_0_out_valid),
    .io_data_0_out_bits(PE_469_io_data_0_out_bits)
  );
  PE PE_470 ( // @[pe.scala 187:13]
    .clock(PE_470_clock),
    .reset(PE_470_reset),
    .io_data_2_out_valid(PE_470_io_data_2_out_valid),
    .io_data_2_out_bits(PE_470_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_470_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_470_io_data_1_in_valid),
    .io_data_1_in_bits(PE_470_io_data_1_in_bits),
    .io_data_1_out_valid(PE_470_io_data_1_out_valid),
    .io_data_1_out_bits(PE_470_io_data_1_out_bits),
    .io_data_0_in_valid(PE_470_io_data_0_in_valid),
    .io_data_0_in_bits(PE_470_io_data_0_in_bits),
    .io_data_0_out_valid(PE_470_io_data_0_out_valid),
    .io_data_0_out_bits(PE_470_io_data_0_out_bits)
  );
  PE PE_471 ( // @[pe.scala 187:13]
    .clock(PE_471_clock),
    .reset(PE_471_reset),
    .io_data_2_out_valid(PE_471_io_data_2_out_valid),
    .io_data_2_out_bits(PE_471_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_471_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_471_io_data_1_in_valid),
    .io_data_1_in_bits(PE_471_io_data_1_in_bits),
    .io_data_1_out_valid(PE_471_io_data_1_out_valid),
    .io_data_1_out_bits(PE_471_io_data_1_out_bits),
    .io_data_0_in_valid(PE_471_io_data_0_in_valid),
    .io_data_0_in_bits(PE_471_io_data_0_in_bits),
    .io_data_0_out_valid(PE_471_io_data_0_out_valid),
    .io_data_0_out_bits(PE_471_io_data_0_out_bits)
  );
  PE PE_472 ( // @[pe.scala 187:13]
    .clock(PE_472_clock),
    .reset(PE_472_reset),
    .io_data_2_out_valid(PE_472_io_data_2_out_valid),
    .io_data_2_out_bits(PE_472_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_472_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_472_io_data_1_in_valid),
    .io_data_1_in_bits(PE_472_io_data_1_in_bits),
    .io_data_1_out_valid(PE_472_io_data_1_out_valid),
    .io_data_1_out_bits(PE_472_io_data_1_out_bits),
    .io_data_0_in_valid(PE_472_io_data_0_in_valid),
    .io_data_0_in_bits(PE_472_io_data_0_in_bits),
    .io_data_0_out_valid(PE_472_io_data_0_out_valid),
    .io_data_0_out_bits(PE_472_io_data_0_out_bits)
  );
  PE PE_473 ( // @[pe.scala 187:13]
    .clock(PE_473_clock),
    .reset(PE_473_reset),
    .io_data_2_out_valid(PE_473_io_data_2_out_valid),
    .io_data_2_out_bits(PE_473_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_473_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_473_io_data_1_in_valid),
    .io_data_1_in_bits(PE_473_io_data_1_in_bits),
    .io_data_1_out_valid(PE_473_io_data_1_out_valid),
    .io_data_1_out_bits(PE_473_io_data_1_out_bits),
    .io_data_0_in_valid(PE_473_io_data_0_in_valid),
    .io_data_0_in_bits(PE_473_io_data_0_in_bits),
    .io_data_0_out_valid(PE_473_io_data_0_out_valid),
    .io_data_0_out_bits(PE_473_io_data_0_out_bits)
  );
  PE PE_474 ( // @[pe.scala 187:13]
    .clock(PE_474_clock),
    .reset(PE_474_reset),
    .io_data_2_out_valid(PE_474_io_data_2_out_valid),
    .io_data_2_out_bits(PE_474_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_474_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_474_io_data_1_in_valid),
    .io_data_1_in_bits(PE_474_io_data_1_in_bits),
    .io_data_1_out_valid(PE_474_io_data_1_out_valid),
    .io_data_1_out_bits(PE_474_io_data_1_out_bits),
    .io_data_0_in_valid(PE_474_io_data_0_in_valid),
    .io_data_0_in_bits(PE_474_io_data_0_in_bits),
    .io_data_0_out_valid(PE_474_io_data_0_out_valid),
    .io_data_0_out_bits(PE_474_io_data_0_out_bits)
  );
  PE PE_475 ( // @[pe.scala 187:13]
    .clock(PE_475_clock),
    .reset(PE_475_reset),
    .io_data_2_out_valid(PE_475_io_data_2_out_valid),
    .io_data_2_out_bits(PE_475_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_475_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_475_io_data_1_in_valid),
    .io_data_1_in_bits(PE_475_io_data_1_in_bits),
    .io_data_1_out_valid(PE_475_io_data_1_out_valid),
    .io_data_1_out_bits(PE_475_io_data_1_out_bits),
    .io_data_0_in_valid(PE_475_io_data_0_in_valid),
    .io_data_0_in_bits(PE_475_io_data_0_in_bits),
    .io_data_0_out_valid(PE_475_io_data_0_out_valid),
    .io_data_0_out_bits(PE_475_io_data_0_out_bits)
  );
  PE PE_476 ( // @[pe.scala 187:13]
    .clock(PE_476_clock),
    .reset(PE_476_reset),
    .io_data_2_out_valid(PE_476_io_data_2_out_valid),
    .io_data_2_out_bits(PE_476_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_476_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_476_io_data_1_in_valid),
    .io_data_1_in_bits(PE_476_io_data_1_in_bits),
    .io_data_1_out_valid(PE_476_io_data_1_out_valid),
    .io_data_1_out_bits(PE_476_io_data_1_out_bits),
    .io_data_0_in_valid(PE_476_io_data_0_in_valid),
    .io_data_0_in_bits(PE_476_io_data_0_in_bits),
    .io_data_0_out_valid(PE_476_io_data_0_out_valid),
    .io_data_0_out_bits(PE_476_io_data_0_out_bits)
  );
  PE PE_477 ( // @[pe.scala 187:13]
    .clock(PE_477_clock),
    .reset(PE_477_reset),
    .io_data_2_out_valid(PE_477_io_data_2_out_valid),
    .io_data_2_out_bits(PE_477_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_477_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_477_io_data_1_in_valid),
    .io_data_1_in_bits(PE_477_io_data_1_in_bits),
    .io_data_1_out_valid(PE_477_io_data_1_out_valid),
    .io_data_1_out_bits(PE_477_io_data_1_out_bits),
    .io_data_0_in_valid(PE_477_io_data_0_in_valid),
    .io_data_0_in_bits(PE_477_io_data_0_in_bits),
    .io_data_0_out_valid(PE_477_io_data_0_out_valid),
    .io_data_0_out_bits(PE_477_io_data_0_out_bits)
  );
  PE PE_478 ( // @[pe.scala 187:13]
    .clock(PE_478_clock),
    .reset(PE_478_reset),
    .io_data_2_out_valid(PE_478_io_data_2_out_valid),
    .io_data_2_out_bits(PE_478_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_478_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_478_io_data_1_in_valid),
    .io_data_1_in_bits(PE_478_io_data_1_in_bits),
    .io_data_1_out_valid(PE_478_io_data_1_out_valid),
    .io_data_1_out_bits(PE_478_io_data_1_out_bits),
    .io_data_0_in_valid(PE_478_io_data_0_in_valid),
    .io_data_0_in_bits(PE_478_io_data_0_in_bits),
    .io_data_0_out_valid(PE_478_io_data_0_out_valid),
    .io_data_0_out_bits(PE_478_io_data_0_out_bits)
  );
  PE PE_479 ( // @[pe.scala 187:13]
    .clock(PE_479_clock),
    .reset(PE_479_reset),
    .io_data_2_out_valid(PE_479_io_data_2_out_valid),
    .io_data_2_out_bits(PE_479_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_479_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_479_io_data_1_in_valid),
    .io_data_1_in_bits(PE_479_io_data_1_in_bits),
    .io_data_1_out_valid(PE_479_io_data_1_out_valid),
    .io_data_1_out_bits(PE_479_io_data_1_out_bits),
    .io_data_0_in_valid(PE_479_io_data_0_in_valid),
    .io_data_0_in_bits(PE_479_io_data_0_in_bits),
    .io_data_0_out_valid(PE_479_io_data_0_out_valid),
    .io_data_0_out_bits(PE_479_io_data_0_out_bits)
  );
  PE PE_480 ( // @[pe.scala 187:13]
    .clock(PE_480_clock),
    .reset(PE_480_reset),
    .io_data_2_out_valid(PE_480_io_data_2_out_valid),
    .io_data_2_out_bits(PE_480_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_480_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_480_io_data_1_in_valid),
    .io_data_1_in_bits(PE_480_io_data_1_in_bits),
    .io_data_1_out_valid(PE_480_io_data_1_out_valid),
    .io_data_1_out_bits(PE_480_io_data_1_out_bits),
    .io_data_0_in_valid(PE_480_io_data_0_in_valid),
    .io_data_0_in_bits(PE_480_io_data_0_in_bits),
    .io_data_0_out_valid(PE_480_io_data_0_out_valid),
    .io_data_0_out_bits(PE_480_io_data_0_out_bits)
  );
  PE PE_481 ( // @[pe.scala 187:13]
    .clock(PE_481_clock),
    .reset(PE_481_reset),
    .io_data_2_out_valid(PE_481_io_data_2_out_valid),
    .io_data_2_out_bits(PE_481_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_481_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_481_io_data_1_in_valid),
    .io_data_1_in_bits(PE_481_io_data_1_in_bits),
    .io_data_1_out_valid(PE_481_io_data_1_out_valid),
    .io_data_1_out_bits(PE_481_io_data_1_out_bits),
    .io_data_0_in_valid(PE_481_io_data_0_in_valid),
    .io_data_0_in_bits(PE_481_io_data_0_in_bits),
    .io_data_0_out_valid(PE_481_io_data_0_out_valid),
    .io_data_0_out_bits(PE_481_io_data_0_out_bits)
  );
  PE PE_482 ( // @[pe.scala 187:13]
    .clock(PE_482_clock),
    .reset(PE_482_reset),
    .io_data_2_out_valid(PE_482_io_data_2_out_valid),
    .io_data_2_out_bits(PE_482_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_482_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_482_io_data_1_in_valid),
    .io_data_1_in_bits(PE_482_io_data_1_in_bits),
    .io_data_1_out_valid(PE_482_io_data_1_out_valid),
    .io_data_1_out_bits(PE_482_io_data_1_out_bits),
    .io_data_0_in_valid(PE_482_io_data_0_in_valid),
    .io_data_0_in_bits(PE_482_io_data_0_in_bits),
    .io_data_0_out_valid(PE_482_io_data_0_out_valid),
    .io_data_0_out_bits(PE_482_io_data_0_out_bits)
  );
  PE PE_483 ( // @[pe.scala 187:13]
    .clock(PE_483_clock),
    .reset(PE_483_reset),
    .io_data_2_out_valid(PE_483_io_data_2_out_valid),
    .io_data_2_out_bits(PE_483_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_483_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_483_io_data_1_in_valid),
    .io_data_1_in_bits(PE_483_io_data_1_in_bits),
    .io_data_1_out_valid(PE_483_io_data_1_out_valid),
    .io_data_1_out_bits(PE_483_io_data_1_out_bits),
    .io_data_0_in_valid(PE_483_io_data_0_in_valid),
    .io_data_0_in_bits(PE_483_io_data_0_in_bits),
    .io_data_0_out_valid(PE_483_io_data_0_out_valid),
    .io_data_0_out_bits(PE_483_io_data_0_out_bits)
  );
  PE PE_484 ( // @[pe.scala 187:13]
    .clock(PE_484_clock),
    .reset(PE_484_reset),
    .io_data_2_out_valid(PE_484_io_data_2_out_valid),
    .io_data_2_out_bits(PE_484_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_484_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_484_io_data_1_in_valid),
    .io_data_1_in_bits(PE_484_io_data_1_in_bits),
    .io_data_1_out_valid(PE_484_io_data_1_out_valid),
    .io_data_1_out_bits(PE_484_io_data_1_out_bits),
    .io_data_0_in_valid(PE_484_io_data_0_in_valid),
    .io_data_0_in_bits(PE_484_io_data_0_in_bits),
    .io_data_0_out_valid(PE_484_io_data_0_out_valid),
    .io_data_0_out_bits(PE_484_io_data_0_out_bits)
  );
  PE PE_485 ( // @[pe.scala 187:13]
    .clock(PE_485_clock),
    .reset(PE_485_reset),
    .io_data_2_out_valid(PE_485_io_data_2_out_valid),
    .io_data_2_out_bits(PE_485_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_485_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_485_io_data_1_in_valid),
    .io_data_1_in_bits(PE_485_io_data_1_in_bits),
    .io_data_1_out_valid(PE_485_io_data_1_out_valid),
    .io_data_1_out_bits(PE_485_io_data_1_out_bits),
    .io_data_0_in_valid(PE_485_io_data_0_in_valid),
    .io_data_0_in_bits(PE_485_io_data_0_in_bits),
    .io_data_0_out_valid(PE_485_io_data_0_out_valid),
    .io_data_0_out_bits(PE_485_io_data_0_out_bits)
  );
  PE PE_486 ( // @[pe.scala 187:13]
    .clock(PE_486_clock),
    .reset(PE_486_reset),
    .io_data_2_out_valid(PE_486_io_data_2_out_valid),
    .io_data_2_out_bits(PE_486_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_486_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_486_io_data_1_in_valid),
    .io_data_1_in_bits(PE_486_io_data_1_in_bits),
    .io_data_1_out_valid(PE_486_io_data_1_out_valid),
    .io_data_1_out_bits(PE_486_io_data_1_out_bits),
    .io_data_0_in_valid(PE_486_io_data_0_in_valid),
    .io_data_0_in_bits(PE_486_io_data_0_in_bits),
    .io_data_0_out_valid(PE_486_io_data_0_out_valid),
    .io_data_0_out_bits(PE_486_io_data_0_out_bits)
  );
  PE PE_487 ( // @[pe.scala 187:13]
    .clock(PE_487_clock),
    .reset(PE_487_reset),
    .io_data_2_out_valid(PE_487_io_data_2_out_valid),
    .io_data_2_out_bits(PE_487_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_487_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_487_io_data_1_in_valid),
    .io_data_1_in_bits(PE_487_io_data_1_in_bits),
    .io_data_1_out_valid(PE_487_io_data_1_out_valid),
    .io_data_1_out_bits(PE_487_io_data_1_out_bits),
    .io_data_0_in_valid(PE_487_io_data_0_in_valid),
    .io_data_0_in_bits(PE_487_io_data_0_in_bits),
    .io_data_0_out_valid(PE_487_io_data_0_out_valid),
    .io_data_0_out_bits(PE_487_io_data_0_out_bits)
  );
  PE PE_488 ( // @[pe.scala 187:13]
    .clock(PE_488_clock),
    .reset(PE_488_reset),
    .io_data_2_out_valid(PE_488_io_data_2_out_valid),
    .io_data_2_out_bits(PE_488_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_488_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_488_io_data_1_in_valid),
    .io_data_1_in_bits(PE_488_io_data_1_in_bits),
    .io_data_1_out_valid(PE_488_io_data_1_out_valid),
    .io_data_1_out_bits(PE_488_io_data_1_out_bits),
    .io_data_0_in_valid(PE_488_io_data_0_in_valid),
    .io_data_0_in_bits(PE_488_io_data_0_in_bits),
    .io_data_0_out_valid(PE_488_io_data_0_out_valid),
    .io_data_0_out_bits(PE_488_io_data_0_out_bits)
  );
  PE PE_489 ( // @[pe.scala 187:13]
    .clock(PE_489_clock),
    .reset(PE_489_reset),
    .io_data_2_out_valid(PE_489_io_data_2_out_valid),
    .io_data_2_out_bits(PE_489_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_489_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_489_io_data_1_in_valid),
    .io_data_1_in_bits(PE_489_io_data_1_in_bits),
    .io_data_1_out_valid(PE_489_io_data_1_out_valid),
    .io_data_1_out_bits(PE_489_io_data_1_out_bits),
    .io_data_0_in_valid(PE_489_io_data_0_in_valid),
    .io_data_0_in_bits(PE_489_io_data_0_in_bits),
    .io_data_0_out_valid(PE_489_io_data_0_out_valid),
    .io_data_0_out_bits(PE_489_io_data_0_out_bits)
  );
  PE PE_490 ( // @[pe.scala 187:13]
    .clock(PE_490_clock),
    .reset(PE_490_reset),
    .io_data_2_out_valid(PE_490_io_data_2_out_valid),
    .io_data_2_out_bits(PE_490_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_490_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_490_io_data_1_in_valid),
    .io_data_1_in_bits(PE_490_io_data_1_in_bits),
    .io_data_1_out_valid(PE_490_io_data_1_out_valid),
    .io_data_1_out_bits(PE_490_io_data_1_out_bits),
    .io_data_0_in_valid(PE_490_io_data_0_in_valid),
    .io_data_0_in_bits(PE_490_io_data_0_in_bits),
    .io_data_0_out_valid(PE_490_io_data_0_out_valid),
    .io_data_0_out_bits(PE_490_io_data_0_out_bits)
  );
  PE PE_491 ( // @[pe.scala 187:13]
    .clock(PE_491_clock),
    .reset(PE_491_reset),
    .io_data_2_out_valid(PE_491_io_data_2_out_valid),
    .io_data_2_out_bits(PE_491_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_491_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_491_io_data_1_in_valid),
    .io_data_1_in_bits(PE_491_io_data_1_in_bits),
    .io_data_1_out_valid(PE_491_io_data_1_out_valid),
    .io_data_1_out_bits(PE_491_io_data_1_out_bits),
    .io_data_0_in_valid(PE_491_io_data_0_in_valid),
    .io_data_0_in_bits(PE_491_io_data_0_in_bits),
    .io_data_0_out_valid(PE_491_io_data_0_out_valid),
    .io_data_0_out_bits(PE_491_io_data_0_out_bits)
  );
  PE PE_492 ( // @[pe.scala 187:13]
    .clock(PE_492_clock),
    .reset(PE_492_reset),
    .io_data_2_out_valid(PE_492_io_data_2_out_valid),
    .io_data_2_out_bits(PE_492_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_492_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_492_io_data_1_in_valid),
    .io_data_1_in_bits(PE_492_io_data_1_in_bits),
    .io_data_1_out_valid(PE_492_io_data_1_out_valid),
    .io_data_1_out_bits(PE_492_io_data_1_out_bits),
    .io_data_0_in_valid(PE_492_io_data_0_in_valid),
    .io_data_0_in_bits(PE_492_io_data_0_in_bits),
    .io_data_0_out_valid(PE_492_io_data_0_out_valid),
    .io_data_0_out_bits(PE_492_io_data_0_out_bits)
  );
  PE PE_493 ( // @[pe.scala 187:13]
    .clock(PE_493_clock),
    .reset(PE_493_reset),
    .io_data_2_out_valid(PE_493_io_data_2_out_valid),
    .io_data_2_out_bits(PE_493_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_493_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_493_io_data_1_in_valid),
    .io_data_1_in_bits(PE_493_io_data_1_in_bits),
    .io_data_1_out_valid(PE_493_io_data_1_out_valid),
    .io_data_1_out_bits(PE_493_io_data_1_out_bits),
    .io_data_0_in_valid(PE_493_io_data_0_in_valid),
    .io_data_0_in_bits(PE_493_io_data_0_in_bits),
    .io_data_0_out_valid(PE_493_io_data_0_out_valid),
    .io_data_0_out_bits(PE_493_io_data_0_out_bits)
  );
  PE PE_494 ( // @[pe.scala 187:13]
    .clock(PE_494_clock),
    .reset(PE_494_reset),
    .io_data_2_out_valid(PE_494_io_data_2_out_valid),
    .io_data_2_out_bits(PE_494_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_494_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_494_io_data_1_in_valid),
    .io_data_1_in_bits(PE_494_io_data_1_in_bits),
    .io_data_1_out_valid(PE_494_io_data_1_out_valid),
    .io_data_1_out_bits(PE_494_io_data_1_out_bits),
    .io_data_0_in_valid(PE_494_io_data_0_in_valid),
    .io_data_0_in_bits(PE_494_io_data_0_in_bits),
    .io_data_0_out_valid(PE_494_io_data_0_out_valid),
    .io_data_0_out_bits(PE_494_io_data_0_out_bits)
  );
  PE PE_495 ( // @[pe.scala 187:13]
    .clock(PE_495_clock),
    .reset(PE_495_reset),
    .io_data_2_out_valid(PE_495_io_data_2_out_valid),
    .io_data_2_out_bits(PE_495_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_495_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_495_io_data_1_in_valid),
    .io_data_1_in_bits(PE_495_io_data_1_in_bits),
    .io_data_1_out_valid(PE_495_io_data_1_out_valid),
    .io_data_1_out_bits(PE_495_io_data_1_out_bits),
    .io_data_0_in_valid(PE_495_io_data_0_in_valid),
    .io_data_0_in_bits(PE_495_io_data_0_in_bits),
    .io_data_0_out_valid(PE_495_io_data_0_out_valid),
    .io_data_0_out_bits(PE_495_io_data_0_out_bits)
  );
  PE PE_496 ( // @[pe.scala 187:13]
    .clock(PE_496_clock),
    .reset(PE_496_reset),
    .io_data_2_out_valid(PE_496_io_data_2_out_valid),
    .io_data_2_out_bits(PE_496_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_496_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_496_io_data_1_in_valid),
    .io_data_1_in_bits(PE_496_io_data_1_in_bits),
    .io_data_1_out_valid(PE_496_io_data_1_out_valid),
    .io_data_1_out_bits(PE_496_io_data_1_out_bits),
    .io_data_0_in_valid(PE_496_io_data_0_in_valid),
    .io_data_0_in_bits(PE_496_io_data_0_in_bits),
    .io_data_0_out_valid(PE_496_io_data_0_out_valid),
    .io_data_0_out_bits(PE_496_io_data_0_out_bits)
  );
  PE PE_497 ( // @[pe.scala 187:13]
    .clock(PE_497_clock),
    .reset(PE_497_reset),
    .io_data_2_out_valid(PE_497_io_data_2_out_valid),
    .io_data_2_out_bits(PE_497_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_497_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_497_io_data_1_in_valid),
    .io_data_1_in_bits(PE_497_io_data_1_in_bits),
    .io_data_1_out_valid(PE_497_io_data_1_out_valid),
    .io_data_1_out_bits(PE_497_io_data_1_out_bits),
    .io_data_0_in_valid(PE_497_io_data_0_in_valid),
    .io_data_0_in_bits(PE_497_io_data_0_in_bits),
    .io_data_0_out_valid(PE_497_io_data_0_out_valid),
    .io_data_0_out_bits(PE_497_io_data_0_out_bits)
  );
  PE PE_498 ( // @[pe.scala 187:13]
    .clock(PE_498_clock),
    .reset(PE_498_reset),
    .io_data_2_out_valid(PE_498_io_data_2_out_valid),
    .io_data_2_out_bits(PE_498_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_498_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_498_io_data_1_in_valid),
    .io_data_1_in_bits(PE_498_io_data_1_in_bits),
    .io_data_1_out_valid(PE_498_io_data_1_out_valid),
    .io_data_1_out_bits(PE_498_io_data_1_out_bits),
    .io_data_0_in_valid(PE_498_io_data_0_in_valid),
    .io_data_0_in_bits(PE_498_io_data_0_in_bits),
    .io_data_0_out_valid(PE_498_io_data_0_out_valid),
    .io_data_0_out_bits(PE_498_io_data_0_out_bits)
  );
  PE PE_499 ( // @[pe.scala 187:13]
    .clock(PE_499_clock),
    .reset(PE_499_reset),
    .io_data_2_out_valid(PE_499_io_data_2_out_valid),
    .io_data_2_out_bits(PE_499_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_499_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_499_io_data_1_in_valid),
    .io_data_1_in_bits(PE_499_io_data_1_in_bits),
    .io_data_1_out_valid(PE_499_io_data_1_out_valid),
    .io_data_1_out_bits(PE_499_io_data_1_out_bits),
    .io_data_0_in_valid(PE_499_io_data_0_in_valid),
    .io_data_0_in_bits(PE_499_io_data_0_in_bits),
    .io_data_0_out_valid(PE_499_io_data_0_out_valid),
    .io_data_0_out_bits(PE_499_io_data_0_out_bits)
  );
  PE PE_500 ( // @[pe.scala 187:13]
    .clock(PE_500_clock),
    .reset(PE_500_reset),
    .io_data_2_out_valid(PE_500_io_data_2_out_valid),
    .io_data_2_out_bits(PE_500_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_500_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_500_io_data_1_in_valid),
    .io_data_1_in_bits(PE_500_io_data_1_in_bits),
    .io_data_1_out_valid(PE_500_io_data_1_out_valid),
    .io_data_1_out_bits(PE_500_io_data_1_out_bits),
    .io_data_0_in_valid(PE_500_io_data_0_in_valid),
    .io_data_0_in_bits(PE_500_io_data_0_in_bits),
    .io_data_0_out_valid(PE_500_io_data_0_out_valid),
    .io_data_0_out_bits(PE_500_io_data_0_out_bits)
  );
  PE PE_501 ( // @[pe.scala 187:13]
    .clock(PE_501_clock),
    .reset(PE_501_reset),
    .io_data_2_out_valid(PE_501_io_data_2_out_valid),
    .io_data_2_out_bits(PE_501_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_501_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_501_io_data_1_in_valid),
    .io_data_1_in_bits(PE_501_io_data_1_in_bits),
    .io_data_1_out_valid(PE_501_io_data_1_out_valid),
    .io_data_1_out_bits(PE_501_io_data_1_out_bits),
    .io_data_0_in_valid(PE_501_io_data_0_in_valid),
    .io_data_0_in_bits(PE_501_io_data_0_in_bits),
    .io_data_0_out_valid(PE_501_io_data_0_out_valid),
    .io_data_0_out_bits(PE_501_io_data_0_out_bits)
  );
  PE PE_502 ( // @[pe.scala 187:13]
    .clock(PE_502_clock),
    .reset(PE_502_reset),
    .io_data_2_out_valid(PE_502_io_data_2_out_valid),
    .io_data_2_out_bits(PE_502_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_502_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_502_io_data_1_in_valid),
    .io_data_1_in_bits(PE_502_io_data_1_in_bits),
    .io_data_1_out_valid(PE_502_io_data_1_out_valid),
    .io_data_1_out_bits(PE_502_io_data_1_out_bits),
    .io_data_0_in_valid(PE_502_io_data_0_in_valid),
    .io_data_0_in_bits(PE_502_io_data_0_in_bits),
    .io_data_0_out_valid(PE_502_io_data_0_out_valid),
    .io_data_0_out_bits(PE_502_io_data_0_out_bits)
  );
  PE PE_503 ( // @[pe.scala 187:13]
    .clock(PE_503_clock),
    .reset(PE_503_reset),
    .io_data_2_out_valid(PE_503_io_data_2_out_valid),
    .io_data_2_out_bits(PE_503_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_503_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_503_io_data_1_in_valid),
    .io_data_1_in_bits(PE_503_io_data_1_in_bits),
    .io_data_1_out_valid(PE_503_io_data_1_out_valid),
    .io_data_1_out_bits(PE_503_io_data_1_out_bits),
    .io_data_0_in_valid(PE_503_io_data_0_in_valid),
    .io_data_0_in_bits(PE_503_io_data_0_in_bits),
    .io_data_0_out_valid(PE_503_io_data_0_out_valid),
    .io_data_0_out_bits(PE_503_io_data_0_out_bits)
  );
  PE PE_504 ( // @[pe.scala 187:13]
    .clock(PE_504_clock),
    .reset(PE_504_reset),
    .io_data_2_out_valid(PE_504_io_data_2_out_valid),
    .io_data_2_out_bits(PE_504_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_504_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_504_io_data_1_in_valid),
    .io_data_1_in_bits(PE_504_io_data_1_in_bits),
    .io_data_1_out_valid(PE_504_io_data_1_out_valid),
    .io_data_1_out_bits(PE_504_io_data_1_out_bits),
    .io_data_0_in_valid(PE_504_io_data_0_in_valid),
    .io_data_0_in_bits(PE_504_io_data_0_in_bits),
    .io_data_0_out_valid(PE_504_io_data_0_out_valid),
    .io_data_0_out_bits(PE_504_io_data_0_out_bits)
  );
  PE PE_505 ( // @[pe.scala 187:13]
    .clock(PE_505_clock),
    .reset(PE_505_reset),
    .io_data_2_out_valid(PE_505_io_data_2_out_valid),
    .io_data_2_out_bits(PE_505_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_505_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_505_io_data_1_in_valid),
    .io_data_1_in_bits(PE_505_io_data_1_in_bits),
    .io_data_1_out_valid(PE_505_io_data_1_out_valid),
    .io_data_1_out_bits(PE_505_io_data_1_out_bits),
    .io_data_0_in_valid(PE_505_io_data_0_in_valid),
    .io_data_0_in_bits(PE_505_io_data_0_in_bits),
    .io_data_0_out_valid(PE_505_io_data_0_out_valid),
    .io_data_0_out_bits(PE_505_io_data_0_out_bits)
  );
  PE PE_506 ( // @[pe.scala 187:13]
    .clock(PE_506_clock),
    .reset(PE_506_reset),
    .io_data_2_out_valid(PE_506_io_data_2_out_valid),
    .io_data_2_out_bits(PE_506_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_506_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_506_io_data_1_in_valid),
    .io_data_1_in_bits(PE_506_io_data_1_in_bits),
    .io_data_1_out_valid(PE_506_io_data_1_out_valid),
    .io_data_1_out_bits(PE_506_io_data_1_out_bits),
    .io_data_0_in_valid(PE_506_io_data_0_in_valid),
    .io_data_0_in_bits(PE_506_io_data_0_in_bits),
    .io_data_0_out_valid(PE_506_io_data_0_out_valid),
    .io_data_0_out_bits(PE_506_io_data_0_out_bits)
  );
  PE PE_507 ( // @[pe.scala 187:13]
    .clock(PE_507_clock),
    .reset(PE_507_reset),
    .io_data_2_out_valid(PE_507_io_data_2_out_valid),
    .io_data_2_out_bits(PE_507_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_507_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_507_io_data_1_in_valid),
    .io_data_1_in_bits(PE_507_io_data_1_in_bits),
    .io_data_1_out_valid(PE_507_io_data_1_out_valid),
    .io_data_1_out_bits(PE_507_io_data_1_out_bits),
    .io_data_0_in_valid(PE_507_io_data_0_in_valid),
    .io_data_0_in_bits(PE_507_io_data_0_in_bits),
    .io_data_0_out_valid(PE_507_io_data_0_out_valid),
    .io_data_0_out_bits(PE_507_io_data_0_out_bits)
  );
  PE PE_508 ( // @[pe.scala 187:13]
    .clock(PE_508_clock),
    .reset(PE_508_reset),
    .io_data_2_out_valid(PE_508_io_data_2_out_valid),
    .io_data_2_out_bits(PE_508_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_508_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_508_io_data_1_in_valid),
    .io_data_1_in_bits(PE_508_io_data_1_in_bits),
    .io_data_1_out_valid(PE_508_io_data_1_out_valid),
    .io_data_1_out_bits(PE_508_io_data_1_out_bits),
    .io_data_0_in_valid(PE_508_io_data_0_in_valid),
    .io_data_0_in_bits(PE_508_io_data_0_in_bits),
    .io_data_0_out_valid(PE_508_io_data_0_out_valid),
    .io_data_0_out_bits(PE_508_io_data_0_out_bits)
  );
  PE PE_509 ( // @[pe.scala 187:13]
    .clock(PE_509_clock),
    .reset(PE_509_reset),
    .io_data_2_out_valid(PE_509_io_data_2_out_valid),
    .io_data_2_out_bits(PE_509_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_509_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_509_io_data_1_in_valid),
    .io_data_1_in_bits(PE_509_io_data_1_in_bits),
    .io_data_1_out_valid(PE_509_io_data_1_out_valid),
    .io_data_1_out_bits(PE_509_io_data_1_out_bits),
    .io_data_0_in_valid(PE_509_io_data_0_in_valid),
    .io_data_0_in_bits(PE_509_io_data_0_in_bits),
    .io_data_0_out_valid(PE_509_io_data_0_out_valid),
    .io_data_0_out_bits(PE_509_io_data_0_out_bits)
  );
  PE PE_510 ( // @[pe.scala 187:13]
    .clock(PE_510_clock),
    .reset(PE_510_reset),
    .io_data_2_out_valid(PE_510_io_data_2_out_valid),
    .io_data_2_out_bits(PE_510_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_510_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_510_io_data_1_in_valid),
    .io_data_1_in_bits(PE_510_io_data_1_in_bits),
    .io_data_1_out_valid(PE_510_io_data_1_out_valid),
    .io_data_1_out_bits(PE_510_io_data_1_out_bits),
    .io_data_0_in_valid(PE_510_io_data_0_in_valid),
    .io_data_0_in_bits(PE_510_io_data_0_in_bits),
    .io_data_0_out_valid(PE_510_io_data_0_out_valid),
    .io_data_0_out_bits(PE_510_io_data_0_out_bits)
  );
  PE PE_511 ( // @[pe.scala 187:13]
    .clock(PE_511_clock),
    .reset(PE_511_reset),
    .io_data_2_out_valid(PE_511_io_data_2_out_valid),
    .io_data_2_out_bits(PE_511_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_511_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_511_io_data_1_in_valid),
    .io_data_1_in_bits(PE_511_io_data_1_in_bits),
    .io_data_1_out_valid(PE_511_io_data_1_out_valid),
    .io_data_1_out_bits(PE_511_io_data_1_out_bits),
    .io_data_0_in_valid(PE_511_io_data_0_in_valid),
    .io_data_0_in_bits(PE_511_io_data_0_in_bits),
    .io_data_0_out_valid(PE_511_io_data_0_out_valid),
    .io_data_0_out_bits(PE_511_io_data_0_out_bits)
  );
  PE PE_512 ( // @[pe.scala 187:13]
    .clock(PE_512_clock),
    .reset(PE_512_reset),
    .io_data_2_out_valid(PE_512_io_data_2_out_valid),
    .io_data_2_out_bits(PE_512_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_512_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_512_io_data_1_in_valid),
    .io_data_1_in_bits(PE_512_io_data_1_in_bits),
    .io_data_1_out_valid(PE_512_io_data_1_out_valid),
    .io_data_1_out_bits(PE_512_io_data_1_out_bits),
    .io_data_0_in_valid(PE_512_io_data_0_in_valid),
    .io_data_0_in_bits(PE_512_io_data_0_in_bits),
    .io_data_0_out_valid(PE_512_io_data_0_out_valid),
    .io_data_0_out_bits(PE_512_io_data_0_out_bits)
  );
  PE PE_513 ( // @[pe.scala 187:13]
    .clock(PE_513_clock),
    .reset(PE_513_reset),
    .io_data_2_out_valid(PE_513_io_data_2_out_valid),
    .io_data_2_out_bits(PE_513_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_513_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_513_io_data_1_in_valid),
    .io_data_1_in_bits(PE_513_io_data_1_in_bits),
    .io_data_1_out_valid(PE_513_io_data_1_out_valid),
    .io_data_1_out_bits(PE_513_io_data_1_out_bits),
    .io_data_0_in_valid(PE_513_io_data_0_in_valid),
    .io_data_0_in_bits(PE_513_io_data_0_in_bits),
    .io_data_0_out_valid(PE_513_io_data_0_out_valid),
    .io_data_0_out_bits(PE_513_io_data_0_out_bits)
  );
  PE PE_514 ( // @[pe.scala 187:13]
    .clock(PE_514_clock),
    .reset(PE_514_reset),
    .io_data_2_out_valid(PE_514_io_data_2_out_valid),
    .io_data_2_out_bits(PE_514_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_514_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_514_io_data_1_in_valid),
    .io_data_1_in_bits(PE_514_io_data_1_in_bits),
    .io_data_1_out_valid(PE_514_io_data_1_out_valid),
    .io_data_1_out_bits(PE_514_io_data_1_out_bits),
    .io_data_0_in_valid(PE_514_io_data_0_in_valid),
    .io_data_0_in_bits(PE_514_io_data_0_in_bits),
    .io_data_0_out_valid(PE_514_io_data_0_out_valid),
    .io_data_0_out_bits(PE_514_io_data_0_out_bits)
  );
  PE PE_515 ( // @[pe.scala 187:13]
    .clock(PE_515_clock),
    .reset(PE_515_reset),
    .io_data_2_out_valid(PE_515_io_data_2_out_valid),
    .io_data_2_out_bits(PE_515_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_515_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_515_io_data_1_in_valid),
    .io_data_1_in_bits(PE_515_io_data_1_in_bits),
    .io_data_1_out_valid(PE_515_io_data_1_out_valid),
    .io_data_1_out_bits(PE_515_io_data_1_out_bits),
    .io_data_0_in_valid(PE_515_io_data_0_in_valid),
    .io_data_0_in_bits(PE_515_io_data_0_in_bits),
    .io_data_0_out_valid(PE_515_io_data_0_out_valid),
    .io_data_0_out_bits(PE_515_io_data_0_out_bits)
  );
  PE PE_516 ( // @[pe.scala 187:13]
    .clock(PE_516_clock),
    .reset(PE_516_reset),
    .io_data_2_out_valid(PE_516_io_data_2_out_valid),
    .io_data_2_out_bits(PE_516_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_516_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_516_io_data_1_in_valid),
    .io_data_1_in_bits(PE_516_io_data_1_in_bits),
    .io_data_1_out_valid(PE_516_io_data_1_out_valid),
    .io_data_1_out_bits(PE_516_io_data_1_out_bits),
    .io_data_0_in_valid(PE_516_io_data_0_in_valid),
    .io_data_0_in_bits(PE_516_io_data_0_in_bits),
    .io_data_0_out_valid(PE_516_io_data_0_out_valid),
    .io_data_0_out_bits(PE_516_io_data_0_out_bits)
  );
  PE PE_517 ( // @[pe.scala 187:13]
    .clock(PE_517_clock),
    .reset(PE_517_reset),
    .io_data_2_out_valid(PE_517_io_data_2_out_valid),
    .io_data_2_out_bits(PE_517_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_517_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_517_io_data_1_in_valid),
    .io_data_1_in_bits(PE_517_io_data_1_in_bits),
    .io_data_1_out_valid(PE_517_io_data_1_out_valid),
    .io_data_1_out_bits(PE_517_io_data_1_out_bits),
    .io_data_0_in_valid(PE_517_io_data_0_in_valid),
    .io_data_0_in_bits(PE_517_io_data_0_in_bits),
    .io_data_0_out_valid(PE_517_io_data_0_out_valid),
    .io_data_0_out_bits(PE_517_io_data_0_out_bits)
  );
  PE PE_518 ( // @[pe.scala 187:13]
    .clock(PE_518_clock),
    .reset(PE_518_reset),
    .io_data_2_out_valid(PE_518_io_data_2_out_valid),
    .io_data_2_out_bits(PE_518_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_518_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_518_io_data_1_in_valid),
    .io_data_1_in_bits(PE_518_io_data_1_in_bits),
    .io_data_1_out_valid(PE_518_io_data_1_out_valid),
    .io_data_1_out_bits(PE_518_io_data_1_out_bits),
    .io_data_0_in_valid(PE_518_io_data_0_in_valid),
    .io_data_0_in_bits(PE_518_io_data_0_in_bits),
    .io_data_0_out_valid(PE_518_io_data_0_out_valid),
    .io_data_0_out_bits(PE_518_io_data_0_out_bits)
  );
  PE PE_519 ( // @[pe.scala 187:13]
    .clock(PE_519_clock),
    .reset(PE_519_reset),
    .io_data_2_out_valid(PE_519_io_data_2_out_valid),
    .io_data_2_out_bits(PE_519_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_519_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_519_io_data_1_in_valid),
    .io_data_1_in_bits(PE_519_io_data_1_in_bits),
    .io_data_1_out_valid(PE_519_io_data_1_out_valid),
    .io_data_1_out_bits(PE_519_io_data_1_out_bits),
    .io_data_0_in_valid(PE_519_io_data_0_in_valid),
    .io_data_0_in_bits(PE_519_io_data_0_in_bits),
    .io_data_0_out_valid(PE_519_io_data_0_out_valid),
    .io_data_0_out_bits(PE_519_io_data_0_out_bits)
  );
  PE PE_520 ( // @[pe.scala 187:13]
    .clock(PE_520_clock),
    .reset(PE_520_reset),
    .io_data_2_out_valid(PE_520_io_data_2_out_valid),
    .io_data_2_out_bits(PE_520_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_520_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_520_io_data_1_in_valid),
    .io_data_1_in_bits(PE_520_io_data_1_in_bits),
    .io_data_1_out_valid(PE_520_io_data_1_out_valid),
    .io_data_1_out_bits(PE_520_io_data_1_out_bits),
    .io_data_0_in_valid(PE_520_io_data_0_in_valid),
    .io_data_0_in_bits(PE_520_io_data_0_in_bits),
    .io_data_0_out_valid(PE_520_io_data_0_out_valid),
    .io_data_0_out_bits(PE_520_io_data_0_out_bits)
  );
  PE PE_521 ( // @[pe.scala 187:13]
    .clock(PE_521_clock),
    .reset(PE_521_reset),
    .io_data_2_out_valid(PE_521_io_data_2_out_valid),
    .io_data_2_out_bits(PE_521_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_521_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_521_io_data_1_in_valid),
    .io_data_1_in_bits(PE_521_io_data_1_in_bits),
    .io_data_1_out_valid(PE_521_io_data_1_out_valid),
    .io_data_1_out_bits(PE_521_io_data_1_out_bits),
    .io_data_0_in_valid(PE_521_io_data_0_in_valid),
    .io_data_0_in_bits(PE_521_io_data_0_in_bits),
    .io_data_0_out_valid(PE_521_io_data_0_out_valid),
    .io_data_0_out_bits(PE_521_io_data_0_out_bits)
  );
  PE PE_522 ( // @[pe.scala 187:13]
    .clock(PE_522_clock),
    .reset(PE_522_reset),
    .io_data_2_out_valid(PE_522_io_data_2_out_valid),
    .io_data_2_out_bits(PE_522_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_522_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_522_io_data_1_in_valid),
    .io_data_1_in_bits(PE_522_io_data_1_in_bits),
    .io_data_1_out_valid(PE_522_io_data_1_out_valid),
    .io_data_1_out_bits(PE_522_io_data_1_out_bits),
    .io_data_0_in_valid(PE_522_io_data_0_in_valid),
    .io_data_0_in_bits(PE_522_io_data_0_in_bits),
    .io_data_0_out_valid(PE_522_io_data_0_out_valid),
    .io_data_0_out_bits(PE_522_io_data_0_out_bits)
  );
  PE PE_523 ( // @[pe.scala 187:13]
    .clock(PE_523_clock),
    .reset(PE_523_reset),
    .io_data_2_out_valid(PE_523_io_data_2_out_valid),
    .io_data_2_out_bits(PE_523_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_523_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_523_io_data_1_in_valid),
    .io_data_1_in_bits(PE_523_io_data_1_in_bits),
    .io_data_1_out_valid(PE_523_io_data_1_out_valid),
    .io_data_1_out_bits(PE_523_io_data_1_out_bits),
    .io_data_0_in_valid(PE_523_io_data_0_in_valid),
    .io_data_0_in_bits(PE_523_io_data_0_in_bits),
    .io_data_0_out_valid(PE_523_io_data_0_out_valid),
    .io_data_0_out_bits(PE_523_io_data_0_out_bits)
  );
  PE PE_524 ( // @[pe.scala 187:13]
    .clock(PE_524_clock),
    .reset(PE_524_reset),
    .io_data_2_out_valid(PE_524_io_data_2_out_valid),
    .io_data_2_out_bits(PE_524_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_524_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_524_io_data_1_in_valid),
    .io_data_1_in_bits(PE_524_io_data_1_in_bits),
    .io_data_1_out_valid(PE_524_io_data_1_out_valid),
    .io_data_1_out_bits(PE_524_io_data_1_out_bits),
    .io_data_0_in_valid(PE_524_io_data_0_in_valid),
    .io_data_0_in_bits(PE_524_io_data_0_in_bits),
    .io_data_0_out_valid(PE_524_io_data_0_out_valid),
    .io_data_0_out_bits(PE_524_io_data_0_out_bits)
  );
  PE PE_525 ( // @[pe.scala 187:13]
    .clock(PE_525_clock),
    .reset(PE_525_reset),
    .io_data_2_out_valid(PE_525_io_data_2_out_valid),
    .io_data_2_out_bits(PE_525_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_525_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_525_io_data_1_in_valid),
    .io_data_1_in_bits(PE_525_io_data_1_in_bits),
    .io_data_1_out_valid(PE_525_io_data_1_out_valid),
    .io_data_1_out_bits(PE_525_io_data_1_out_bits),
    .io_data_0_in_valid(PE_525_io_data_0_in_valid),
    .io_data_0_in_bits(PE_525_io_data_0_in_bits),
    .io_data_0_out_valid(PE_525_io_data_0_out_valid),
    .io_data_0_out_bits(PE_525_io_data_0_out_bits)
  );
  PE PE_526 ( // @[pe.scala 187:13]
    .clock(PE_526_clock),
    .reset(PE_526_reset),
    .io_data_2_out_valid(PE_526_io_data_2_out_valid),
    .io_data_2_out_bits(PE_526_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_526_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_526_io_data_1_in_valid),
    .io_data_1_in_bits(PE_526_io_data_1_in_bits),
    .io_data_1_out_valid(PE_526_io_data_1_out_valid),
    .io_data_1_out_bits(PE_526_io_data_1_out_bits),
    .io_data_0_in_valid(PE_526_io_data_0_in_valid),
    .io_data_0_in_bits(PE_526_io_data_0_in_bits),
    .io_data_0_out_valid(PE_526_io_data_0_out_valid),
    .io_data_0_out_bits(PE_526_io_data_0_out_bits)
  );
  PE PE_527 ( // @[pe.scala 187:13]
    .clock(PE_527_clock),
    .reset(PE_527_reset),
    .io_data_2_out_valid(PE_527_io_data_2_out_valid),
    .io_data_2_out_bits(PE_527_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_527_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_527_io_data_1_in_valid),
    .io_data_1_in_bits(PE_527_io_data_1_in_bits),
    .io_data_1_out_valid(PE_527_io_data_1_out_valid),
    .io_data_1_out_bits(PE_527_io_data_1_out_bits),
    .io_data_0_in_valid(PE_527_io_data_0_in_valid),
    .io_data_0_in_bits(PE_527_io_data_0_in_bits),
    .io_data_0_out_valid(PE_527_io_data_0_out_valid),
    .io_data_0_out_bits(PE_527_io_data_0_out_bits)
  );
  PE PE_528 ( // @[pe.scala 187:13]
    .clock(PE_528_clock),
    .reset(PE_528_reset),
    .io_data_2_out_valid(PE_528_io_data_2_out_valid),
    .io_data_2_out_bits(PE_528_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_528_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_528_io_data_1_in_valid),
    .io_data_1_in_bits(PE_528_io_data_1_in_bits),
    .io_data_1_out_valid(PE_528_io_data_1_out_valid),
    .io_data_1_out_bits(PE_528_io_data_1_out_bits),
    .io_data_0_in_valid(PE_528_io_data_0_in_valid),
    .io_data_0_in_bits(PE_528_io_data_0_in_bits),
    .io_data_0_out_valid(PE_528_io_data_0_out_valid),
    .io_data_0_out_bits(PE_528_io_data_0_out_bits)
  );
  PE PE_529 ( // @[pe.scala 187:13]
    .clock(PE_529_clock),
    .reset(PE_529_reset),
    .io_data_2_out_valid(PE_529_io_data_2_out_valid),
    .io_data_2_out_bits(PE_529_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_529_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_529_io_data_1_in_valid),
    .io_data_1_in_bits(PE_529_io_data_1_in_bits),
    .io_data_1_out_valid(PE_529_io_data_1_out_valid),
    .io_data_1_out_bits(PE_529_io_data_1_out_bits),
    .io_data_0_in_valid(PE_529_io_data_0_in_valid),
    .io_data_0_in_bits(PE_529_io_data_0_in_bits),
    .io_data_0_out_valid(PE_529_io_data_0_out_valid),
    .io_data_0_out_bits(PE_529_io_data_0_out_bits)
  );
  PE PE_530 ( // @[pe.scala 187:13]
    .clock(PE_530_clock),
    .reset(PE_530_reset),
    .io_data_2_out_valid(PE_530_io_data_2_out_valid),
    .io_data_2_out_bits(PE_530_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_530_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_530_io_data_1_in_valid),
    .io_data_1_in_bits(PE_530_io_data_1_in_bits),
    .io_data_1_out_valid(PE_530_io_data_1_out_valid),
    .io_data_1_out_bits(PE_530_io_data_1_out_bits),
    .io_data_0_in_valid(PE_530_io_data_0_in_valid),
    .io_data_0_in_bits(PE_530_io_data_0_in_bits),
    .io_data_0_out_valid(PE_530_io_data_0_out_valid),
    .io_data_0_out_bits(PE_530_io_data_0_out_bits)
  );
  PE PE_531 ( // @[pe.scala 187:13]
    .clock(PE_531_clock),
    .reset(PE_531_reset),
    .io_data_2_out_valid(PE_531_io_data_2_out_valid),
    .io_data_2_out_bits(PE_531_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_531_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_531_io_data_1_in_valid),
    .io_data_1_in_bits(PE_531_io_data_1_in_bits),
    .io_data_1_out_valid(PE_531_io_data_1_out_valid),
    .io_data_1_out_bits(PE_531_io_data_1_out_bits),
    .io_data_0_in_valid(PE_531_io_data_0_in_valid),
    .io_data_0_in_bits(PE_531_io_data_0_in_bits),
    .io_data_0_out_valid(PE_531_io_data_0_out_valid),
    .io_data_0_out_bits(PE_531_io_data_0_out_bits)
  );
  PE PE_532 ( // @[pe.scala 187:13]
    .clock(PE_532_clock),
    .reset(PE_532_reset),
    .io_data_2_out_valid(PE_532_io_data_2_out_valid),
    .io_data_2_out_bits(PE_532_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_532_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_532_io_data_1_in_valid),
    .io_data_1_in_bits(PE_532_io_data_1_in_bits),
    .io_data_1_out_valid(PE_532_io_data_1_out_valid),
    .io_data_1_out_bits(PE_532_io_data_1_out_bits),
    .io_data_0_in_valid(PE_532_io_data_0_in_valid),
    .io_data_0_in_bits(PE_532_io_data_0_in_bits),
    .io_data_0_out_valid(PE_532_io_data_0_out_valid),
    .io_data_0_out_bits(PE_532_io_data_0_out_bits)
  );
  PE PE_533 ( // @[pe.scala 187:13]
    .clock(PE_533_clock),
    .reset(PE_533_reset),
    .io_data_2_out_valid(PE_533_io_data_2_out_valid),
    .io_data_2_out_bits(PE_533_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_533_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_533_io_data_1_in_valid),
    .io_data_1_in_bits(PE_533_io_data_1_in_bits),
    .io_data_1_out_valid(PE_533_io_data_1_out_valid),
    .io_data_1_out_bits(PE_533_io_data_1_out_bits),
    .io_data_0_in_valid(PE_533_io_data_0_in_valid),
    .io_data_0_in_bits(PE_533_io_data_0_in_bits),
    .io_data_0_out_valid(PE_533_io_data_0_out_valid),
    .io_data_0_out_bits(PE_533_io_data_0_out_bits)
  );
  PE PE_534 ( // @[pe.scala 187:13]
    .clock(PE_534_clock),
    .reset(PE_534_reset),
    .io_data_2_out_valid(PE_534_io_data_2_out_valid),
    .io_data_2_out_bits(PE_534_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_534_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_534_io_data_1_in_valid),
    .io_data_1_in_bits(PE_534_io_data_1_in_bits),
    .io_data_1_out_valid(PE_534_io_data_1_out_valid),
    .io_data_1_out_bits(PE_534_io_data_1_out_bits),
    .io_data_0_in_valid(PE_534_io_data_0_in_valid),
    .io_data_0_in_bits(PE_534_io_data_0_in_bits),
    .io_data_0_out_valid(PE_534_io_data_0_out_valid),
    .io_data_0_out_bits(PE_534_io_data_0_out_bits)
  );
  PE PE_535 ( // @[pe.scala 187:13]
    .clock(PE_535_clock),
    .reset(PE_535_reset),
    .io_data_2_out_valid(PE_535_io_data_2_out_valid),
    .io_data_2_out_bits(PE_535_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_535_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_535_io_data_1_in_valid),
    .io_data_1_in_bits(PE_535_io_data_1_in_bits),
    .io_data_1_out_valid(PE_535_io_data_1_out_valid),
    .io_data_1_out_bits(PE_535_io_data_1_out_bits),
    .io_data_0_in_valid(PE_535_io_data_0_in_valid),
    .io_data_0_in_bits(PE_535_io_data_0_in_bits),
    .io_data_0_out_valid(PE_535_io_data_0_out_valid),
    .io_data_0_out_bits(PE_535_io_data_0_out_bits)
  );
  PE PE_536 ( // @[pe.scala 187:13]
    .clock(PE_536_clock),
    .reset(PE_536_reset),
    .io_data_2_out_valid(PE_536_io_data_2_out_valid),
    .io_data_2_out_bits(PE_536_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_536_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_536_io_data_1_in_valid),
    .io_data_1_in_bits(PE_536_io_data_1_in_bits),
    .io_data_1_out_valid(PE_536_io_data_1_out_valid),
    .io_data_1_out_bits(PE_536_io_data_1_out_bits),
    .io_data_0_in_valid(PE_536_io_data_0_in_valid),
    .io_data_0_in_bits(PE_536_io_data_0_in_bits),
    .io_data_0_out_valid(PE_536_io_data_0_out_valid),
    .io_data_0_out_bits(PE_536_io_data_0_out_bits)
  );
  PE PE_537 ( // @[pe.scala 187:13]
    .clock(PE_537_clock),
    .reset(PE_537_reset),
    .io_data_2_out_valid(PE_537_io_data_2_out_valid),
    .io_data_2_out_bits(PE_537_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_537_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_537_io_data_1_in_valid),
    .io_data_1_in_bits(PE_537_io_data_1_in_bits),
    .io_data_1_out_valid(PE_537_io_data_1_out_valid),
    .io_data_1_out_bits(PE_537_io_data_1_out_bits),
    .io_data_0_in_valid(PE_537_io_data_0_in_valid),
    .io_data_0_in_bits(PE_537_io_data_0_in_bits),
    .io_data_0_out_valid(PE_537_io_data_0_out_valid),
    .io_data_0_out_bits(PE_537_io_data_0_out_bits)
  );
  PE PE_538 ( // @[pe.scala 187:13]
    .clock(PE_538_clock),
    .reset(PE_538_reset),
    .io_data_2_out_valid(PE_538_io_data_2_out_valid),
    .io_data_2_out_bits(PE_538_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_538_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_538_io_data_1_in_valid),
    .io_data_1_in_bits(PE_538_io_data_1_in_bits),
    .io_data_1_out_valid(PE_538_io_data_1_out_valid),
    .io_data_1_out_bits(PE_538_io_data_1_out_bits),
    .io_data_0_in_valid(PE_538_io_data_0_in_valid),
    .io_data_0_in_bits(PE_538_io_data_0_in_bits),
    .io_data_0_out_valid(PE_538_io_data_0_out_valid),
    .io_data_0_out_bits(PE_538_io_data_0_out_bits)
  );
  PE PE_539 ( // @[pe.scala 187:13]
    .clock(PE_539_clock),
    .reset(PE_539_reset),
    .io_data_2_out_valid(PE_539_io_data_2_out_valid),
    .io_data_2_out_bits(PE_539_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_539_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_539_io_data_1_in_valid),
    .io_data_1_in_bits(PE_539_io_data_1_in_bits),
    .io_data_1_out_valid(PE_539_io_data_1_out_valid),
    .io_data_1_out_bits(PE_539_io_data_1_out_bits),
    .io_data_0_in_valid(PE_539_io_data_0_in_valid),
    .io_data_0_in_bits(PE_539_io_data_0_in_bits),
    .io_data_0_out_valid(PE_539_io_data_0_out_valid),
    .io_data_0_out_bits(PE_539_io_data_0_out_bits)
  );
  PE PE_540 ( // @[pe.scala 187:13]
    .clock(PE_540_clock),
    .reset(PE_540_reset),
    .io_data_2_out_valid(PE_540_io_data_2_out_valid),
    .io_data_2_out_bits(PE_540_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_540_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_540_io_data_1_in_valid),
    .io_data_1_in_bits(PE_540_io_data_1_in_bits),
    .io_data_1_out_valid(PE_540_io_data_1_out_valid),
    .io_data_1_out_bits(PE_540_io_data_1_out_bits),
    .io_data_0_in_valid(PE_540_io_data_0_in_valid),
    .io_data_0_in_bits(PE_540_io_data_0_in_bits),
    .io_data_0_out_valid(PE_540_io_data_0_out_valid),
    .io_data_0_out_bits(PE_540_io_data_0_out_bits)
  );
  PE PE_541 ( // @[pe.scala 187:13]
    .clock(PE_541_clock),
    .reset(PE_541_reset),
    .io_data_2_out_valid(PE_541_io_data_2_out_valid),
    .io_data_2_out_bits(PE_541_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_541_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_541_io_data_1_in_valid),
    .io_data_1_in_bits(PE_541_io_data_1_in_bits),
    .io_data_1_out_valid(PE_541_io_data_1_out_valid),
    .io_data_1_out_bits(PE_541_io_data_1_out_bits),
    .io_data_0_in_valid(PE_541_io_data_0_in_valid),
    .io_data_0_in_bits(PE_541_io_data_0_in_bits),
    .io_data_0_out_valid(PE_541_io_data_0_out_valid),
    .io_data_0_out_bits(PE_541_io_data_0_out_bits)
  );
  PE PE_542 ( // @[pe.scala 187:13]
    .clock(PE_542_clock),
    .reset(PE_542_reset),
    .io_data_2_out_valid(PE_542_io_data_2_out_valid),
    .io_data_2_out_bits(PE_542_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_542_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_542_io_data_1_in_valid),
    .io_data_1_in_bits(PE_542_io_data_1_in_bits),
    .io_data_1_out_valid(PE_542_io_data_1_out_valid),
    .io_data_1_out_bits(PE_542_io_data_1_out_bits),
    .io_data_0_in_valid(PE_542_io_data_0_in_valid),
    .io_data_0_in_bits(PE_542_io_data_0_in_bits),
    .io_data_0_out_valid(PE_542_io_data_0_out_valid),
    .io_data_0_out_bits(PE_542_io_data_0_out_bits)
  );
  PE PE_543 ( // @[pe.scala 187:13]
    .clock(PE_543_clock),
    .reset(PE_543_reset),
    .io_data_2_out_valid(PE_543_io_data_2_out_valid),
    .io_data_2_out_bits(PE_543_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_543_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_543_io_data_1_in_valid),
    .io_data_1_in_bits(PE_543_io_data_1_in_bits),
    .io_data_1_out_valid(PE_543_io_data_1_out_valid),
    .io_data_1_out_bits(PE_543_io_data_1_out_bits),
    .io_data_0_in_valid(PE_543_io_data_0_in_valid),
    .io_data_0_in_bits(PE_543_io_data_0_in_bits),
    .io_data_0_out_valid(PE_543_io_data_0_out_valid),
    .io_data_0_out_bits(PE_543_io_data_0_out_bits)
  );
  PE PE_544 ( // @[pe.scala 187:13]
    .clock(PE_544_clock),
    .reset(PE_544_reset),
    .io_data_2_out_valid(PE_544_io_data_2_out_valid),
    .io_data_2_out_bits(PE_544_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_544_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_544_io_data_1_in_valid),
    .io_data_1_in_bits(PE_544_io_data_1_in_bits),
    .io_data_1_out_valid(PE_544_io_data_1_out_valid),
    .io_data_1_out_bits(PE_544_io_data_1_out_bits),
    .io_data_0_in_valid(PE_544_io_data_0_in_valid),
    .io_data_0_in_bits(PE_544_io_data_0_in_bits),
    .io_data_0_out_valid(PE_544_io_data_0_out_valid),
    .io_data_0_out_bits(PE_544_io_data_0_out_bits)
  );
  PE PE_545 ( // @[pe.scala 187:13]
    .clock(PE_545_clock),
    .reset(PE_545_reset),
    .io_data_2_out_valid(PE_545_io_data_2_out_valid),
    .io_data_2_out_bits(PE_545_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_545_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_545_io_data_1_in_valid),
    .io_data_1_in_bits(PE_545_io_data_1_in_bits),
    .io_data_1_out_valid(PE_545_io_data_1_out_valid),
    .io_data_1_out_bits(PE_545_io_data_1_out_bits),
    .io_data_0_in_valid(PE_545_io_data_0_in_valid),
    .io_data_0_in_bits(PE_545_io_data_0_in_bits),
    .io_data_0_out_valid(PE_545_io_data_0_out_valid),
    .io_data_0_out_bits(PE_545_io_data_0_out_bits)
  );
  PE PE_546 ( // @[pe.scala 187:13]
    .clock(PE_546_clock),
    .reset(PE_546_reset),
    .io_data_2_out_valid(PE_546_io_data_2_out_valid),
    .io_data_2_out_bits(PE_546_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_546_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_546_io_data_1_in_valid),
    .io_data_1_in_bits(PE_546_io_data_1_in_bits),
    .io_data_1_out_valid(PE_546_io_data_1_out_valid),
    .io_data_1_out_bits(PE_546_io_data_1_out_bits),
    .io_data_0_in_valid(PE_546_io_data_0_in_valid),
    .io_data_0_in_bits(PE_546_io_data_0_in_bits),
    .io_data_0_out_valid(PE_546_io_data_0_out_valid),
    .io_data_0_out_bits(PE_546_io_data_0_out_bits)
  );
  PE PE_547 ( // @[pe.scala 187:13]
    .clock(PE_547_clock),
    .reset(PE_547_reset),
    .io_data_2_out_valid(PE_547_io_data_2_out_valid),
    .io_data_2_out_bits(PE_547_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_547_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_547_io_data_1_in_valid),
    .io_data_1_in_bits(PE_547_io_data_1_in_bits),
    .io_data_1_out_valid(PE_547_io_data_1_out_valid),
    .io_data_1_out_bits(PE_547_io_data_1_out_bits),
    .io_data_0_in_valid(PE_547_io_data_0_in_valid),
    .io_data_0_in_bits(PE_547_io_data_0_in_bits),
    .io_data_0_out_valid(PE_547_io_data_0_out_valid),
    .io_data_0_out_bits(PE_547_io_data_0_out_bits)
  );
  PE PE_548 ( // @[pe.scala 187:13]
    .clock(PE_548_clock),
    .reset(PE_548_reset),
    .io_data_2_out_valid(PE_548_io_data_2_out_valid),
    .io_data_2_out_bits(PE_548_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_548_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_548_io_data_1_in_valid),
    .io_data_1_in_bits(PE_548_io_data_1_in_bits),
    .io_data_1_out_valid(PE_548_io_data_1_out_valid),
    .io_data_1_out_bits(PE_548_io_data_1_out_bits),
    .io_data_0_in_valid(PE_548_io_data_0_in_valid),
    .io_data_0_in_bits(PE_548_io_data_0_in_bits),
    .io_data_0_out_valid(PE_548_io_data_0_out_valid),
    .io_data_0_out_bits(PE_548_io_data_0_out_bits)
  );
  PE PE_549 ( // @[pe.scala 187:13]
    .clock(PE_549_clock),
    .reset(PE_549_reset),
    .io_data_2_out_valid(PE_549_io_data_2_out_valid),
    .io_data_2_out_bits(PE_549_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_549_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_549_io_data_1_in_valid),
    .io_data_1_in_bits(PE_549_io_data_1_in_bits),
    .io_data_1_out_valid(PE_549_io_data_1_out_valid),
    .io_data_1_out_bits(PE_549_io_data_1_out_bits),
    .io_data_0_in_valid(PE_549_io_data_0_in_valid),
    .io_data_0_in_bits(PE_549_io_data_0_in_bits),
    .io_data_0_out_valid(PE_549_io_data_0_out_valid),
    .io_data_0_out_bits(PE_549_io_data_0_out_bits)
  );
  PE PE_550 ( // @[pe.scala 187:13]
    .clock(PE_550_clock),
    .reset(PE_550_reset),
    .io_data_2_out_valid(PE_550_io_data_2_out_valid),
    .io_data_2_out_bits(PE_550_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_550_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_550_io_data_1_in_valid),
    .io_data_1_in_bits(PE_550_io_data_1_in_bits),
    .io_data_1_out_valid(PE_550_io_data_1_out_valid),
    .io_data_1_out_bits(PE_550_io_data_1_out_bits),
    .io_data_0_in_valid(PE_550_io_data_0_in_valid),
    .io_data_0_in_bits(PE_550_io_data_0_in_bits),
    .io_data_0_out_valid(PE_550_io_data_0_out_valid),
    .io_data_0_out_bits(PE_550_io_data_0_out_bits)
  );
  PE PE_551 ( // @[pe.scala 187:13]
    .clock(PE_551_clock),
    .reset(PE_551_reset),
    .io_data_2_out_valid(PE_551_io_data_2_out_valid),
    .io_data_2_out_bits(PE_551_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_551_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_551_io_data_1_in_valid),
    .io_data_1_in_bits(PE_551_io_data_1_in_bits),
    .io_data_1_out_valid(PE_551_io_data_1_out_valid),
    .io_data_1_out_bits(PE_551_io_data_1_out_bits),
    .io_data_0_in_valid(PE_551_io_data_0_in_valid),
    .io_data_0_in_bits(PE_551_io_data_0_in_bits),
    .io_data_0_out_valid(PE_551_io_data_0_out_valid),
    .io_data_0_out_bits(PE_551_io_data_0_out_bits)
  );
  PE PE_552 ( // @[pe.scala 187:13]
    .clock(PE_552_clock),
    .reset(PE_552_reset),
    .io_data_2_out_valid(PE_552_io_data_2_out_valid),
    .io_data_2_out_bits(PE_552_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_552_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_552_io_data_1_in_valid),
    .io_data_1_in_bits(PE_552_io_data_1_in_bits),
    .io_data_1_out_valid(PE_552_io_data_1_out_valid),
    .io_data_1_out_bits(PE_552_io_data_1_out_bits),
    .io_data_0_in_valid(PE_552_io_data_0_in_valid),
    .io_data_0_in_bits(PE_552_io_data_0_in_bits),
    .io_data_0_out_valid(PE_552_io_data_0_out_valid),
    .io_data_0_out_bits(PE_552_io_data_0_out_bits)
  );
  PE PE_553 ( // @[pe.scala 187:13]
    .clock(PE_553_clock),
    .reset(PE_553_reset),
    .io_data_2_out_valid(PE_553_io_data_2_out_valid),
    .io_data_2_out_bits(PE_553_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_553_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_553_io_data_1_in_valid),
    .io_data_1_in_bits(PE_553_io_data_1_in_bits),
    .io_data_1_out_valid(PE_553_io_data_1_out_valid),
    .io_data_1_out_bits(PE_553_io_data_1_out_bits),
    .io_data_0_in_valid(PE_553_io_data_0_in_valid),
    .io_data_0_in_bits(PE_553_io_data_0_in_bits),
    .io_data_0_out_valid(PE_553_io_data_0_out_valid),
    .io_data_0_out_bits(PE_553_io_data_0_out_bits)
  );
  PE PE_554 ( // @[pe.scala 187:13]
    .clock(PE_554_clock),
    .reset(PE_554_reset),
    .io_data_2_out_valid(PE_554_io_data_2_out_valid),
    .io_data_2_out_bits(PE_554_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_554_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_554_io_data_1_in_valid),
    .io_data_1_in_bits(PE_554_io_data_1_in_bits),
    .io_data_1_out_valid(PE_554_io_data_1_out_valid),
    .io_data_1_out_bits(PE_554_io_data_1_out_bits),
    .io_data_0_in_valid(PE_554_io_data_0_in_valid),
    .io_data_0_in_bits(PE_554_io_data_0_in_bits),
    .io_data_0_out_valid(PE_554_io_data_0_out_valid),
    .io_data_0_out_bits(PE_554_io_data_0_out_bits)
  );
  PE PE_555 ( // @[pe.scala 187:13]
    .clock(PE_555_clock),
    .reset(PE_555_reset),
    .io_data_2_out_valid(PE_555_io_data_2_out_valid),
    .io_data_2_out_bits(PE_555_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_555_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_555_io_data_1_in_valid),
    .io_data_1_in_bits(PE_555_io_data_1_in_bits),
    .io_data_1_out_valid(PE_555_io_data_1_out_valid),
    .io_data_1_out_bits(PE_555_io_data_1_out_bits),
    .io_data_0_in_valid(PE_555_io_data_0_in_valid),
    .io_data_0_in_bits(PE_555_io_data_0_in_bits),
    .io_data_0_out_valid(PE_555_io_data_0_out_valid),
    .io_data_0_out_bits(PE_555_io_data_0_out_bits)
  );
  PE PE_556 ( // @[pe.scala 187:13]
    .clock(PE_556_clock),
    .reset(PE_556_reset),
    .io_data_2_out_valid(PE_556_io_data_2_out_valid),
    .io_data_2_out_bits(PE_556_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_556_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_556_io_data_1_in_valid),
    .io_data_1_in_bits(PE_556_io_data_1_in_bits),
    .io_data_1_out_valid(PE_556_io_data_1_out_valid),
    .io_data_1_out_bits(PE_556_io_data_1_out_bits),
    .io_data_0_in_valid(PE_556_io_data_0_in_valid),
    .io_data_0_in_bits(PE_556_io_data_0_in_bits),
    .io_data_0_out_valid(PE_556_io_data_0_out_valid),
    .io_data_0_out_bits(PE_556_io_data_0_out_bits)
  );
  PE PE_557 ( // @[pe.scala 187:13]
    .clock(PE_557_clock),
    .reset(PE_557_reset),
    .io_data_2_out_valid(PE_557_io_data_2_out_valid),
    .io_data_2_out_bits(PE_557_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_557_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_557_io_data_1_in_valid),
    .io_data_1_in_bits(PE_557_io_data_1_in_bits),
    .io_data_1_out_valid(PE_557_io_data_1_out_valid),
    .io_data_1_out_bits(PE_557_io_data_1_out_bits),
    .io_data_0_in_valid(PE_557_io_data_0_in_valid),
    .io_data_0_in_bits(PE_557_io_data_0_in_bits),
    .io_data_0_out_valid(PE_557_io_data_0_out_valid),
    .io_data_0_out_bits(PE_557_io_data_0_out_bits)
  );
  PE PE_558 ( // @[pe.scala 187:13]
    .clock(PE_558_clock),
    .reset(PE_558_reset),
    .io_data_2_out_valid(PE_558_io_data_2_out_valid),
    .io_data_2_out_bits(PE_558_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_558_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_558_io_data_1_in_valid),
    .io_data_1_in_bits(PE_558_io_data_1_in_bits),
    .io_data_1_out_valid(PE_558_io_data_1_out_valid),
    .io_data_1_out_bits(PE_558_io_data_1_out_bits),
    .io_data_0_in_valid(PE_558_io_data_0_in_valid),
    .io_data_0_in_bits(PE_558_io_data_0_in_bits),
    .io_data_0_out_valid(PE_558_io_data_0_out_valid),
    .io_data_0_out_bits(PE_558_io_data_0_out_bits)
  );
  PE PE_559 ( // @[pe.scala 187:13]
    .clock(PE_559_clock),
    .reset(PE_559_reset),
    .io_data_2_out_valid(PE_559_io_data_2_out_valid),
    .io_data_2_out_bits(PE_559_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_559_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_559_io_data_1_in_valid),
    .io_data_1_in_bits(PE_559_io_data_1_in_bits),
    .io_data_1_out_valid(PE_559_io_data_1_out_valid),
    .io_data_1_out_bits(PE_559_io_data_1_out_bits),
    .io_data_0_in_valid(PE_559_io_data_0_in_valid),
    .io_data_0_in_bits(PE_559_io_data_0_in_bits),
    .io_data_0_out_valid(PE_559_io_data_0_out_valid),
    .io_data_0_out_bits(PE_559_io_data_0_out_bits)
  );
  PE PE_560 ( // @[pe.scala 187:13]
    .clock(PE_560_clock),
    .reset(PE_560_reset),
    .io_data_2_out_valid(PE_560_io_data_2_out_valid),
    .io_data_2_out_bits(PE_560_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_560_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_560_io_data_1_in_valid),
    .io_data_1_in_bits(PE_560_io_data_1_in_bits),
    .io_data_1_out_valid(PE_560_io_data_1_out_valid),
    .io_data_1_out_bits(PE_560_io_data_1_out_bits),
    .io_data_0_in_valid(PE_560_io_data_0_in_valid),
    .io_data_0_in_bits(PE_560_io_data_0_in_bits),
    .io_data_0_out_valid(PE_560_io_data_0_out_valid),
    .io_data_0_out_bits(PE_560_io_data_0_out_bits)
  );
  PE PE_561 ( // @[pe.scala 187:13]
    .clock(PE_561_clock),
    .reset(PE_561_reset),
    .io_data_2_out_valid(PE_561_io_data_2_out_valid),
    .io_data_2_out_bits(PE_561_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_561_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_561_io_data_1_in_valid),
    .io_data_1_in_bits(PE_561_io_data_1_in_bits),
    .io_data_1_out_valid(PE_561_io_data_1_out_valid),
    .io_data_1_out_bits(PE_561_io_data_1_out_bits),
    .io_data_0_in_valid(PE_561_io_data_0_in_valid),
    .io_data_0_in_bits(PE_561_io_data_0_in_bits),
    .io_data_0_out_valid(PE_561_io_data_0_out_valid),
    .io_data_0_out_bits(PE_561_io_data_0_out_bits)
  );
  PE PE_562 ( // @[pe.scala 187:13]
    .clock(PE_562_clock),
    .reset(PE_562_reset),
    .io_data_2_out_valid(PE_562_io_data_2_out_valid),
    .io_data_2_out_bits(PE_562_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_562_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_562_io_data_1_in_valid),
    .io_data_1_in_bits(PE_562_io_data_1_in_bits),
    .io_data_1_out_valid(PE_562_io_data_1_out_valid),
    .io_data_1_out_bits(PE_562_io_data_1_out_bits),
    .io_data_0_in_valid(PE_562_io_data_0_in_valid),
    .io_data_0_in_bits(PE_562_io_data_0_in_bits),
    .io_data_0_out_valid(PE_562_io_data_0_out_valid),
    .io_data_0_out_bits(PE_562_io_data_0_out_bits)
  );
  PE PE_563 ( // @[pe.scala 187:13]
    .clock(PE_563_clock),
    .reset(PE_563_reset),
    .io_data_2_out_valid(PE_563_io_data_2_out_valid),
    .io_data_2_out_bits(PE_563_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_563_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_563_io_data_1_in_valid),
    .io_data_1_in_bits(PE_563_io_data_1_in_bits),
    .io_data_1_out_valid(PE_563_io_data_1_out_valid),
    .io_data_1_out_bits(PE_563_io_data_1_out_bits),
    .io_data_0_in_valid(PE_563_io_data_0_in_valid),
    .io_data_0_in_bits(PE_563_io_data_0_in_bits),
    .io_data_0_out_valid(PE_563_io_data_0_out_valid),
    .io_data_0_out_bits(PE_563_io_data_0_out_bits)
  );
  PE PE_564 ( // @[pe.scala 187:13]
    .clock(PE_564_clock),
    .reset(PE_564_reset),
    .io_data_2_out_valid(PE_564_io_data_2_out_valid),
    .io_data_2_out_bits(PE_564_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_564_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_564_io_data_1_in_valid),
    .io_data_1_in_bits(PE_564_io_data_1_in_bits),
    .io_data_1_out_valid(PE_564_io_data_1_out_valid),
    .io_data_1_out_bits(PE_564_io_data_1_out_bits),
    .io_data_0_in_valid(PE_564_io_data_0_in_valid),
    .io_data_0_in_bits(PE_564_io_data_0_in_bits),
    .io_data_0_out_valid(PE_564_io_data_0_out_valid),
    .io_data_0_out_bits(PE_564_io_data_0_out_bits)
  );
  PE PE_565 ( // @[pe.scala 187:13]
    .clock(PE_565_clock),
    .reset(PE_565_reset),
    .io_data_2_out_valid(PE_565_io_data_2_out_valid),
    .io_data_2_out_bits(PE_565_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_565_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_565_io_data_1_in_valid),
    .io_data_1_in_bits(PE_565_io_data_1_in_bits),
    .io_data_1_out_valid(PE_565_io_data_1_out_valid),
    .io_data_1_out_bits(PE_565_io_data_1_out_bits),
    .io_data_0_in_valid(PE_565_io_data_0_in_valid),
    .io_data_0_in_bits(PE_565_io_data_0_in_bits),
    .io_data_0_out_valid(PE_565_io_data_0_out_valid),
    .io_data_0_out_bits(PE_565_io_data_0_out_bits)
  );
  PE PE_566 ( // @[pe.scala 187:13]
    .clock(PE_566_clock),
    .reset(PE_566_reset),
    .io_data_2_out_valid(PE_566_io_data_2_out_valid),
    .io_data_2_out_bits(PE_566_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_566_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_566_io_data_1_in_valid),
    .io_data_1_in_bits(PE_566_io_data_1_in_bits),
    .io_data_1_out_valid(PE_566_io_data_1_out_valid),
    .io_data_1_out_bits(PE_566_io_data_1_out_bits),
    .io_data_0_in_valid(PE_566_io_data_0_in_valid),
    .io_data_0_in_bits(PE_566_io_data_0_in_bits),
    .io_data_0_out_valid(PE_566_io_data_0_out_valid),
    .io_data_0_out_bits(PE_566_io_data_0_out_bits)
  );
  PE PE_567 ( // @[pe.scala 187:13]
    .clock(PE_567_clock),
    .reset(PE_567_reset),
    .io_data_2_out_valid(PE_567_io_data_2_out_valid),
    .io_data_2_out_bits(PE_567_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_567_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_567_io_data_1_in_valid),
    .io_data_1_in_bits(PE_567_io_data_1_in_bits),
    .io_data_1_out_valid(PE_567_io_data_1_out_valid),
    .io_data_1_out_bits(PE_567_io_data_1_out_bits),
    .io_data_0_in_valid(PE_567_io_data_0_in_valid),
    .io_data_0_in_bits(PE_567_io_data_0_in_bits),
    .io_data_0_out_valid(PE_567_io_data_0_out_valid),
    .io_data_0_out_bits(PE_567_io_data_0_out_bits)
  );
  PE PE_568 ( // @[pe.scala 187:13]
    .clock(PE_568_clock),
    .reset(PE_568_reset),
    .io_data_2_out_valid(PE_568_io_data_2_out_valid),
    .io_data_2_out_bits(PE_568_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_568_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_568_io_data_1_in_valid),
    .io_data_1_in_bits(PE_568_io_data_1_in_bits),
    .io_data_1_out_valid(PE_568_io_data_1_out_valid),
    .io_data_1_out_bits(PE_568_io_data_1_out_bits),
    .io_data_0_in_valid(PE_568_io_data_0_in_valid),
    .io_data_0_in_bits(PE_568_io_data_0_in_bits),
    .io_data_0_out_valid(PE_568_io_data_0_out_valid),
    .io_data_0_out_bits(PE_568_io_data_0_out_bits)
  );
  PE PE_569 ( // @[pe.scala 187:13]
    .clock(PE_569_clock),
    .reset(PE_569_reset),
    .io_data_2_out_valid(PE_569_io_data_2_out_valid),
    .io_data_2_out_bits(PE_569_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_569_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_569_io_data_1_in_valid),
    .io_data_1_in_bits(PE_569_io_data_1_in_bits),
    .io_data_1_out_valid(PE_569_io_data_1_out_valid),
    .io_data_1_out_bits(PE_569_io_data_1_out_bits),
    .io_data_0_in_valid(PE_569_io_data_0_in_valid),
    .io_data_0_in_bits(PE_569_io_data_0_in_bits),
    .io_data_0_out_valid(PE_569_io_data_0_out_valid),
    .io_data_0_out_bits(PE_569_io_data_0_out_bits)
  );
  PE PE_570 ( // @[pe.scala 187:13]
    .clock(PE_570_clock),
    .reset(PE_570_reset),
    .io_data_2_out_valid(PE_570_io_data_2_out_valid),
    .io_data_2_out_bits(PE_570_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_570_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_570_io_data_1_in_valid),
    .io_data_1_in_bits(PE_570_io_data_1_in_bits),
    .io_data_1_out_valid(PE_570_io_data_1_out_valid),
    .io_data_1_out_bits(PE_570_io_data_1_out_bits),
    .io_data_0_in_valid(PE_570_io_data_0_in_valid),
    .io_data_0_in_bits(PE_570_io_data_0_in_bits),
    .io_data_0_out_valid(PE_570_io_data_0_out_valid),
    .io_data_0_out_bits(PE_570_io_data_0_out_bits)
  );
  PE PE_571 ( // @[pe.scala 187:13]
    .clock(PE_571_clock),
    .reset(PE_571_reset),
    .io_data_2_out_valid(PE_571_io_data_2_out_valid),
    .io_data_2_out_bits(PE_571_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_571_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_571_io_data_1_in_valid),
    .io_data_1_in_bits(PE_571_io_data_1_in_bits),
    .io_data_1_out_valid(PE_571_io_data_1_out_valid),
    .io_data_1_out_bits(PE_571_io_data_1_out_bits),
    .io_data_0_in_valid(PE_571_io_data_0_in_valid),
    .io_data_0_in_bits(PE_571_io_data_0_in_bits),
    .io_data_0_out_valid(PE_571_io_data_0_out_valid),
    .io_data_0_out_bits(PE_571_io_data_0_out_bits)
  );
  PE PE_572 ( // @[pe.scala 187:13]
    .clock(PE_572_clock),
    .reset(PE_572_reset),
    .io_data_2_out_valid(PE_572_io_data_2_out_valid),
    .io_data_2_out_bits(PE_572_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_572_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_572_io_data_1_in_valid),
    .io_data_1_in_bits(PE_572_io_data_1_in_bits),
    .io_data_1_out_valid(PE_572_io_data_1_out_valid),
    .io_data_1_out_bits(PE_572_io_data_1_out_bits),
    .io_data_0_in_valid(PE_572_io_data_0_in_valid),
    .io_data_0_in_bits(PE_572_io_data_0_in_bits),
    .io_data_0_out_valid(PE_572_io_data_0_out_valid),
    .io_data_0_out_bits(PE_572_io_data_0_out_bits)
  );
  PE PE_573 ( // @[pe.scala 187:13]
    .clock(PE_573_clock),
    .reset(PE_573_reset),
    .io_data_2_out_valid(PE_573_io_data_2_out_valid),
    .io_data_2_out_bits(PE_573_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_573_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_573_io_data_1_in_valid),
    .io_data_1_in_bits(PE_573_io_data_1_in_bits),
    .io_data_1_out_valid(PE_573_io_data_1_out_valid),
    .io_data_1_out_bits(PE_573_io_data_1_out_bits),
    .io_data_0_in_valid(PE_573_io_data_0_in_valid),
    .io_data_0_in_bits(PE_573_io_data_0_in_bits),
    .io_data_0_out_valid(PE_573_io_data_0_out_valid),
    .io_data_0_out_bits(PE_573_io_data_0_out_bits)
  );
  PE PE_574 ( // @[pe.scala 187:13]
    .clock(PE_574_clock),
    .reset(PE_574_reset),
    .io_data_2_out_valid(PE_574_io_data_2_out_valid),
    .io_data_2_out_bits(PE_574_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_574_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_574_io_data_1_in_valid),
    .io_data_1_in_bits(PE_574_io_data_1_in_bits),
    .io_data_1_out_valid(PE_574_io_data_1_out_valid),
    .io_data_1_out_bits(PE_574_io_data_1_out_bits),
    .io_data_0_in_valid(PE_574_io_data_0_in_valid),
    .io_data_0_in_bits(PE_574_io_data_0_in_bits),
    .io_data_0_out_valid(PE_574_io_data_0_out_valid),
    .io_data_0_out_bits(PE_574_io_data_0_out_bits)
  );
  PE PE_575 ( // @[pe.scala 187:13]
    .clock(PE_575_clock),
    .reset(PE_575_reset),
    .io_data_2_out_valid(PE_575_io_data_2_out_valid),
    .io_data_2_out_bits(PE_575_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_575_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_575_io_data_1_in_valid),
    .io_data_1_in_bits(PE_575_io_data_1_in_bits),
    .io_data_1_out_valid(PE_575_io_data_1_out_valid),
    .io_data_1_out_bits(PE_575_io_data_1_out_bits),
    .io_data_0_in_valid(PE_575_io_data_0_in_valid),
    .io_data_0_in_bits(PE_575_io_data_0_in_bits),
    .io_data_0_out_valid(PE_575_io_data_0_out_valid),
    .io_data_0_out_bits(PE_575_io_data_0_out_bits)
  );
  PE PE_576 ( // @[pe.scala 187:13]
    .clock(PE_576_clock),
    .reset(PE_576_reset),
    .io_data_2_out_valid(PE_576_io_data_2_out_valid),
    .io_data_2_out_bits(PE_576_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_576_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_576_io_data_1_in_valid),
    .io_data_1_in_bits(PE_576_io_data_1_in_bits),
    .io_data_1_out_valid(PE_576_io_data_1_out_valid),
    .io_data_1_out_bits(PE_576_io_data_1_out_bits),
    .io_data_0_in_valid(PE_576_io_data_0_in_valid),
    .io_data_0_in_bits(PE_576_io_data_0_in_bits),
    .io_data_0_out_valid(PE_576_io_data_0_out_valid),
    .io_data_0_out_bits(PE_576_io_data_0_out_bits)
  );
  PE PE_577 ( // @[pe.scala 187:13]
    .clock(PE_577_clock),
    .reset(PE_577_reset),
    .io_data_2_out_valid(PE_577_io_data_2_out_valid),
    .io_data_2_out_bits(PE_577_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_577_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_577_io_data_1_in_valid),
    .io_data_1_in_bits(PE_577_io_data_1_in_bits),
    .io_data_1_out_valid(PE_577_io_data_1_out_valid),
    .io_data_1_out_bits(PE_577_io_data_1_out_bits),
    .io_data_0_in_valid(PE_577_io_data_0_in_valid),
    .io_data_0_in_bits(PE_577_io_data_0_in_bits),
    .io_data_0_out_valid(PE_577_io_data_0_out_valid),
    .io_data_0_out_bits(PE_577_io_data_0_out_bits)
  );
  PE PE_578 ( // @[pe.scala 187:13]
    .clock(PE_578_clock),
    .reset(PE_578_reset),
    .io_data_2_out_valid(PE_578_io_data_2_out_valid),
    .io_data_2_out_bits(PE_578_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_578_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_578_io_data_1_in_valid),
    .io_data_1_in_bits(PE_578_io_data_1_in_bits),
    .io_data_1_out_valid(PE_578_io_data_1_out_valid),
    .io_data_1_out_bits(PE_578_io_data_1_out_bits),
    .io_data_0_in_valid(PE_578_io_data_0_in_valid),
    .io_data_0_in_bits(PE_578_io_data_0_in_bits),
    .io_data_0_out_valid(PE_578_io_data_0_out_valid),
    .io_data_0_out_bits(PE_578_io_data_0_out_bits)
  );
  PE PE_579 ( // @[pe.scala 187:13]
    .clock(PE_579_clock),
    .reset(PE_579_reset),
    .io_data_2_out_valid(PE_579_io_data_2_out_valid),
    .io_data_2_out_bits(PE_579_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_579_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_579_io_data_1_in_valid),
    .io_data_1_in_bits(PE_579_io_data_1_in_bits),
    .io_data_1_out_valid(PE_579_io_data_1_out_valid),
    .io_data_1_out_bits(PE_579_io_data_1_out_bits),
    .io_data_0_in_valid(PE_579_io_data_0_in_valid),
    .io_data_0_in_bits(PE_579_io_data_0_in_bits),
    .io_data_0_out_valid(PE_579_io_data_0_out_valid),
    .io_data_0_out_bits(PE_579_io_data_0_out_bits)
  );
  PE PE_580 ( // @[pe.scala 187:13]
    .clock(PE_580_clock),
    .reset(PE_580_reset),
    .io_data_2_out_valid(PE_580_io_data_2_out_valid),
    .io_data_2_out_bits(PE_580_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_580_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_580_io_data_1_in_valid),
    .io_data_1_in_bits(PE_580_io_data_1_in_bits),
    .io_data_1_out_valid(PE_580_io_data_1_out_valid),
    .io_data_1_out_bits(PE_580_io_data_1_out_bits),
    .io_data_0_in_valid(PE_580_io_data_0_in_valid),
    .io_data_0_in_bits(PE_580_io_data_0_in_bits),
    .io_data_0_out_valid(PE_580_io_data_0_out_valid),
    .io_data_0_out_bits(PE_580_io_data_0_out_bits)
  );
  PE PE_581 ( // @[pe.scala 187:13]
    .clock(PE_581_clock),
    .reset(PE_581_reset),
    .io_data_2_out_valid(PE_581_io_data_2_out_valid),
    .io_data_2_out_bits(PE_581_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_581_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_581_io_data_1_in_valid),
    .io_data_1_in_bits(PE_581_io_data_1_in_bits),
    .io_data_1_out_valid(PE_581_io_data_1_out_valid),
    .io_data_1_out_bits(PE_581_io_data_1_out_bits),
    .io_data_0_in_valid(PE_581_io_data_0_in_valid),
    .io_data_0_in_bits(PE_581_io_data_0_in_bits),
    .io_data_0_out_valid(PE_581_io_data_0_out_valid),
    .io_data_0_out_bits(PE_581_io_data_0_out_bits)
  );
  PE PE_582 ( // @[pe.scala 187:13]
    .clock(PE_582_clock),
    .reset(PE_582_reset),
    .io_data_2_out_valid(PE_582_io_data_2_out_valid),
    .io_data_2_out_bits(PE_582_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_582_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_582_io_data_1_in_valid),
    .io_data_1_in_bits(PE_582_io_data_1_in_bits),
    .io_data_1_out_valid(PE_582_io_data_1_out_valid),
    .io_data_1_out_bits(PE_582_io_data_1_out_bits),
    .io_data_0_in_valid(PE_582_io_data_0_in_valid),
    .io_data_0_in_bits(PE_582_io_data_0_in_bits),
    .io_data_0_out_valid(PE_582_io_data_0_out_valid),
    .io_data_0_out_bits(PE_582_io_data_0_out_bits)
  );
  PE PE_583 ( // @[pe.scala 187:13]
    .clock(PE_583_clock),
    .reset(PE_583_reset),
    .io_data_2_out_valid(PE_583_io_data_2_out_valid),
    .io_data_2_out_bits(PE_583_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_583_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_583_io_data_1_in_valid),
    .io_data_1_in_bits(PE_583_io_data_1_in_bits),
    .io_data_1_out_valid(PE_583_io_data_1_out_valid),
    .io_data_1_out_bits(PE_583_io_data_1_out_bits),
    .io_data_0_in_valid(PE_583_io_data_0_in_valid),
    .io_data_0_in_bits(PE_583_io_data_0_in_bits),
    .io_data_0_out_valid(PE_583_io_data_0_out_valid),
    .io_data_0_out_bits(PE_583_io_data_0_out_bits)
  );
  PE PE_584 ( // @[pe.scala 187:13]
    .clock(PE_584_clock),
    .reset(PE_584_reset),
    .io_data_2_out_valid(PE_584_io_data_2_out_valid),
    .io_data_2_out_bits(PE_584_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_584_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_584_io_data_1_in_valid),
    .io_data_1_in_bits(PE_584_io_data_1_in_bits),
    .io_data_1_out_valid(PE_584_io_data_1_out_valid),
    .io_data_1_out_bits(PE_584_io_data_1_out_bits),
    .io_data_0_in_valid(PE_584_io_data_0_in_valid),
    .io_data_0_in_bits(PE_584_io_data_0_in_bits),
    .io_data_0_out_valid(PE_584_io_data_0_out_valid),
    .io_data_0_out_bits(PE_584_io_data_0_out_bits)
  );
  PE PE_585 ( // @[pe.scala 187:13]
    .clock(PE_585_clock),
    .reset(PE_585_reset),
    .io_data_2_out_valid(PE_585_io_data_2_out_valid),
    .io_data_2_out_bits(PE_585_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_585_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_585_io_data_1_in_valid),
    .io_data_1_in_bits(PE_585_io_data_1_in_bits),
    .io_data_1_out_valid(PE_585_io_data_1_out_valid),
    .io_data_1_out_bits(PE_585_io_data_1_out_bits),
    .io_data_0_in_valid(PE_585_io_data_0_in_valid),
    .io_data_0_in_bits(PE_585_io_data_0_in_bits),
    .io_data_0_out_valid(PE_585_io_data_0_out_valid),
    .io_data_0_out_bits(PE_585_io_data_0_out_bits)
  );
  PE PE_586 ( // @[pe.scala 187:13]
    .clock(PE_586_clock),
    .reset(PE_586_reset),
    .io_data_2_out_valid(PE_586_io_data_2_out_valid),
    .io_data_2_out_bits(PE_586_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_586_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_586_io_data_1_in_valid),
    .io_data_1_in_bits(PE_586_io_data_1_in_bits),
    .io_data_1_out_valid(PE_586_io_data_1_out_valid),
    .io_data_1_out_bits(PE_586_io_data_1_out_bits),
    .io_data_0_in_valid(PE_586_io_data_0_in_valid),
    .io_data_0_in_bits(PE_586_io_data_0_in_bits),
    .io_data_0_out_valid(PE_586_io_data_0_out_valid),
    .io_data_0_out_bits(PE_586_io_data_0_out_bits)
  );
  PE PE_587 ( // @[pe.scala 187:13]
    .clock(PE_587_clock),
    .reset(PE_587_reset),
    .io_data_2_out_valid(PE_587_io_data_2_out_valid),
    .io_data_2_out_bits(PE_587_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_587_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_587_io_data_1_in_valid),
    .io_data_1_in_bits(PE_587_io_data_1_in_bits),
    .io_data_1_out_valid(PE_587_io_data_1_out_valid),
    .io_data_1_out_bits(PE_587_io_data_1_out_bits),
    .io_data_0_in_valid(PE_587_io_data_0_in_valid),
    .io_data_0_in_bits(PE_587_io_data_0_in_bits),
    .io_data_0_out_valid(PE_587_io_data_0_out_valid),
    .io_data_0_out_bits(PE_587_io_data_0_out_bits)
  );
  PE PE_588 ( // @[pe.scala 187:13]
    .clock(PE_588_clock),
    .reset(PE_588_reset),
    .io_data_2_out_valid(PE_588_io_data_2_out_valid),
    .io_data_2_out_bits(PE_588_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_588_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_588_io_data_1_in_valid),
    .io_data_1_in_bits(PE_588_io_data_1_in_bits),
    .io_data_1_out_valid(PE_588_io_data_1_out_valid),
    .io_data_1_out_bits(PE_588_io_data_1_out_bits),
    .io_data_0_in_valid(PE_588_io_data_0_in_valid),
    .io_data_0_in_bits(PE_588_io_data_0_in_bits),
    .io_data_0_out_valid(PE_588_io_data_0_out_valid),
    .io_data_0_out_bits(PE_588_io_data_0_out_bits)
  );
  PE PE_589 ( // @[pe.scala 187:13]
    .clock(PE_589_clock),
    .reset(PE_589_reset),
    .io_data_2_out_valid(PE_589_io_data_2_out_valid),
    .io_data_2_out_bits(PE_589_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_589_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_589_io_data_1_in_valid),
    .io_data_1_in_bits(PE_589_io_data_1_in_bits),
    .io_data_1_out_valid(PE_589_io_data_1_out_valid),
    .io_data_1_out_bits(PE_589_io_data_1_out_bits),
    .io_data_0_in_valid(PE_589_io_data_0_in_valid),
    .io_data_0_in_bits(PE_589_io_data_0_in_bits),
    .io_data_0_out_valid(PE_589_io_data_0_out_valid),
    .io_data_0_out_bits(PE_589_io_data_0_out_bits)
  );
  PE PE_590 ( // @[pe.scala 187:13]
    .clock(PE_590_clock),
    .reset(PE_590_reset),
    .io_data_2_out_valid(PE_590_io_data_2_out_valid),
    .io_data_2_out_bits(PE_590_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_590_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_590_io_data_1_in_valid),
    .io_data_1_in_bits(PE_590_io_data_1_in_bits),
    .io_data_1_out_valid(PE_590_io_data_1_out_valid),
    .io_data_1_out_bits(PE_590_io_data_1_out_bits),
    .io_data_0_in_valid(PE_590_io_data_0_in_valid),
    .io_data_0_in_bits(PE_590_io_data_0_in_bits),
    .io_data_0_out_valid(PE_590_io_data_0_out_valid),
    .io_data_0_out_bits(PE_590_io_data_0_out_bits)
  );
  PE PE_591 ( // @[pe.scala 187:13]
    .clock(PE_591_clock),
    .reset(PE_591_reset),
    .io_data_2_out_valid(PE_591_io_data_2_out_valid),
    .io_data_2_out_bits(PE_591_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_591_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_591_io_data_1_in_valid),
    .io_data_1_in_bits(PE_591_io_data_1_in_bits),
    .io_data_1_out_valid(PE_591_io_data_1_out_valid),
    .io_data_1_out_bits(PE_591_io_data_1_out_bits),
    .io_data_0_in_valid(PE_591_io_data_0_in_valid),
    .io_data_0_in_bits(PE_591_io_data_0_in_bits),
    .io_data_0_out_valid(PE_591_io_data_0_out_valid),
    .io_data_0_out_bits(PE_591_io_data_0_out_bits)
  );
  PE PE_592 ( // @[pe.scala 187:13]
    .clock(PE_592_clock),
    .reset(PE_592_reset),
    .io_data_2_out_valid(PE_592_io_data_2_out_valid),
    .io_data_2_out_bits(PE_592_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_592_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_592_io_data_1_in_valid),
    .io_data_1_in_bits(PE_592_io_data_1_in_bits),
    .io_data_1_out_valid(PE_592_io_data_1_out_valid),
    .io_data_1_out_bits(PE_592_io_data_1_out_bits),
    .io_data_0_in_valid(PE_592_io_data_0_in_valid),
    .io_data_0_in_bits(PE_592_io_data_0_in_bits),
    .io_data_0_out_valid(PE_592_io_data_0_out_valid),
    .io_data_0_out_bits(PE_592_io_data_0_out_bits)
  );
  PE PE_593 ( // @[pe.scala 187:13]
    .clock(PE_593_clock),
    .reset(PE_593_reset),
    .io_data_2_out_valid(PE_593_io_data_2_out_valid),
    .io_data_2_out_bits(PE_593_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_593_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_593_io_data_1_in_valid),
    .io_data_1_in_bits(PE_593_io_data_1_in_bits),
    .io_data_1_out_valid(PE_593_io_data_1_out_valid),
    .io_data_1_out_bits(PE_593_io_data_1_out_bits),
    .io_data_0_in_valid(PE_593_io_data_0_in_valid),
    .io_data_0_in_bits(PE_593_io_data_0_in_bits),
    .io_data_0_out_valid(PE_593_io_data_0_out_valid),
    .io_data_0_out_bits(PE_593_io_data_0_out_bits)
  );
  PE PE_594 ( // @[pe.scala 187:13]
    .clock(PE_594_clock),
    .reset(PE_594_reset),
    .io_data_2_out_valid(PE_594_io_data_2_out_valid),
    .io_data_2_out_bits(PE_594_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_594_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_594_io_data_1_in_valid),
    .io_data_1_in_bits(PE_594_io_data_1_in_bits),
    .io_data_1_out_valid(PE_594_io_data_1_out_valid),
    .io_data_1_out_bits(PE_594_io_data_1_out_bits),
    .io_data_0_in_valid(PE_594_io_data_0_in_valid),
    .io_data_0_in_bits(PE_594_io_data_0_in_bits),
    .io_data_0_out_valid(PE_594_io_data_0_out_valid),
    .io_data_0_out_bits(PE_594_io_data_0_out_bits)
  );
  PE PE_595 ( // @[pe.scala 187:13]
    .clock(PE_595_clock),
    .reset(PE_595_reset),
    .io_data_2_out_valid(PE_595_io_data_2_out_valid),
    .io_data_2_out_bits(PE_595_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_595_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_595_io_data_1_in_valid),
    .io_data_1_in_bits(PE_595_io_data_1_in_bits),
    .io_data_1_out_valid(PE_595_io_data_1_out_valid),
    .io_data_1_out_bits(PE_595_io_data_1_out_bits),
    .io_data_0_in_valid(PE_595_io_data_0_in_valid),
    .io_data_0_in_bits(PE_595_io_data_0_in_bits),
    .io_data_0_out_valid(PE_595_io_data_0_out_valid),
    .io_data_0_out_bits(PE_595_io_data_0_out_bits)
  );
  PE PE_596 ( // @[pe.scala 187:13]
    .clock(PE_596_clock),
    .reset(PE_596_reset),
    .io_data_2_out_valid(PE_596_io_data_2_out_valid),
    .io_data_2_out_bits(PE_596_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_596_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_596_io_data_1_in_valid),
    .io_data_1_in_bits(PE_596_io_data_1_in_bits),
    .io_data_1_out_valid(PE_596_io_data_1_out_valid),
    .io_data_1_out_bits(PE_596_io_data_1_out_bits),
    .io_data_0_in_valid(PE_596_io_data_0_in_valid),
    .io_data_0_in_bits(PE_596_io_data_0_in_bits),
    .io_data_0_out_valid(PE_596_io_data_0_out_valid),
    .io_data_0_out_bits(PE_596_io_data_0_out_bits)
  );
  PE PE_597 ( // @[pe.scala 187:13]
    .clock(PE_597_clock),
    .reset(PE_597_reset),
    .io_data_2_out_valid(PE_597_io_data_2_out_valid),
    .io_data_2_out_bits(PE_597_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_597_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_597_io_data_1_in_valid),
    .io_data_1_in_bits(PE_597_io_data_1_in_bits),
    .io_data_1_out_valid(PE_597_io_data_1_out_valid),
    .io_data_1_out_bits(PE_597_io_data_1_out_bits),
    .io_data_0_in_valid(PE_597_io_data_0_in_valid),
    .io_data_0_in_bits(PE_597_io_data_0_in_bits),
    .io_data_0_out_valid(PE_597_io_data_0_out_valid),
    .io_data_0_out_bits(PE_597_io_data_0_out_bits)
  );
  PE PE_598 ( // @[pe.scala 187:13]
    .clock(PE_598_clock),
    .reset(PE_598_reset),
    .io_data_2_out_valid(PE_598_io_data_2_out_valid),
    .io_data_2_out_bits(PE_598_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_598_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_598_io_data_1_in_valid),
    .io_data_1_in_bits(PE_598_io_data_1_in_bits),
    .io_data_1_out_valid(PE_598_io_data_1_out_valid),
    .io_data_1_out_bits(PE_598_io_data_1_out_bits),
    .io_data_0_in_valid(PE_598_io_data_0_in_valid),
    .io_data_0_in_bits(PE_598_io_data_0_in_bits),
    .io_data_0_out_valid(PE_598_io_data_0_out_valid),
    .io_data_0_out_bits(PE_598_io_data_0_out_bits)
  );
  PE PE_599 ( // @[pe.scala 187:13]
    .clock(PE_599_clock),
    .reset(PE_599_reset),
    .io_data_2_out_valid(PE_599_io_data_2_out_valid),
    .io_data_2_out_bits(PE_599_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_599_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_599_io_data_1_in_valid),
    .io_data_1_in_bits(PE_599_io_data_1_in_bits),
    .io_data_1_out_valid(PE_599_io_data_1_out_valid),
    .io_data_1_out_bits(PE_599_io_data_1_out_bits),
    .io_data_0_in_valid(PE_599_io_data_0_in_valid),
    .io_data_0_in_bits(PE_599_io_data_0_in_bits),
    .io_data_0_out_valid(PE_599_io_data_0_out_valid),
    .io_data_0_out_bits(PE_599_io_data_0_out_bits)
  );
  PE PE_600 ( // @[pe.scala 187:13]
    .clock(PE_600_clock),
    .reset(PE_600_reset),
    .io_data_2_out_valid(PE_600_io_data_2_out_valid),
    .io_data_2_out_bits(PE_600_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_600_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_600_io_data_1_in_valid),
    .io_data_1_in_bits(PE_600_io_data_1_in_bits),
    .io_data_1_out_valid(PE_600_io_data_1_out_valid),
    .io_data_1_out_bits(PE_600_io_data_1_out_bits),
    .io_data_0_in_valid(PE_600_io_data_0_in_valid),
    .io_data_0_in_bits(PE_600_io_data_0_in_bits),
    .io_data_0_out_valid(PE_600_io_data_0_out_valid),
    .io_data_0_out_bits(PE_600_io_data_0_out_bits)
  );
  PE PE_601 ( // @[pe.scala 187:13]
    .clock(PE_601_clock),
    .reset(PE_601_reset),
    .io_data_2_out_valid(PE_601_io_data_2_out_valid),
    .io_data_2_out_bits(PE_601_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_601_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_601_io_data_1_in_valid),
    .io_data_1_in_bits(PE_601_io_data_1_in_bits),
    .io_data_1_out_valid(PE_601_io_data_1_out_valid),
    .io_data_1_out_bits(PE_601_io_data_1_out_bits),
    .io_data_0_in_valid(PE_601_io_data_0_in_valid),
    .io_data_0_in_bits(PE_601_io_data_0_in_bits),
    .io_data_0_out_valid(PE_601_io_data_0_out_valid),
    .io_data_0_out_bits(PE_601_io_data_0_out_bits)
  );
  PE PE_602 ( // @[pe.scala 187:13]
    .clock(PE_602_clock),
    .reset(PE_602_reset),
    .io_data_2_out_valid(PE_602_io_data_2_out_valid),
    .io_data_2_out_bits(PE_602_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_602_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_602_io_data_1_in_valid),
    .io_data_1_in_bits(PE_602_io_data_1_in_bits),
    .io_data_1_out_valid(PE_602_io_data_1_out_valid),
    .io_data_1_out_bits(PE_602_io_data_1_out_bits),
    .io_data_0_in_valid(PE_602_io_data_0_in_valid),
    .io_data_0_in_bits(PE_602_io_data_0_in_bits),
    .io_data_0_out_valid(PE_602_io_data_0_out_valid),
    .io_data_0_out_bits(PE_602_io_data_0_out_bits)
  );
  PE PE_603 ( // @[pe.scala 187:13]
    .clock(PE_603_clock),
    .reset(PE_603_reset),
    .io_data_2_out_valid(PE_603_io_data_2_out_valid),
    .io_data_2_out_bits(PE_603_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_603_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_603_io_data_1_in_valid),
    .io_data_1_in_bits(PE_603_io_data_1_in_bits),
    .io_data_1_out_valid(PE_603_io_data_1_out_valid),
    .io_data_1_out_bits(PE_603_io_data_1_out_bits),
    .io_data_0_in_valid(PE_603_io_data_0_in_valid),
    .io_data_0_in_bits(PE_603_io_data_0_in_bits),
    .io_data_0_out_valid(PE_603_io_data_0_out_valid),
    .io_data_0_out_bits(PE_603_io_data_0_out_bits)
  );
  PE PE_604 ( // @[pe.scala 187:13]
    .clock(PE_604_clock),
    .reset(PE_604_reset),
    .io_data_2_out_valid(PE_604_io_data_2_out_valid),
    .io_data_2_out_bits(PE_604_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_604_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_604_io_data_1_in_valid),
    .io_data_1_in_bits(PE_604_io_data_1_in_bits),
    .io_data_1_out_valid(PE_604_io_data_1_out_valid),
    .io_data_1_out_bits(PE_604_io_data_1_out_bits),
    .io_data_0_in_valid(PE_604_io_data_0_in_valid),
    .io_data_0_in_bits(PE_604_io_data_0_in_bits),
    .io_data_0_out_valid(PE_604_io_data_0_out_valid),
    .io_data_0_out_bits(PE_604_io_data_0_out_bits)
  );
  PE PE_605 ( // @[pe.scala 187:13]
    .clock(PE_605_clock),
    .reset(PE_605_reset),
    .io_data_2_out_valid(PE_605_io_data_2_out_valid),
    .io_data_2_out_bits(PE_605_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_605_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_605_io_data_1_in_valid),
    .io_data_1_in_bits(PE_605_io_data_1_in_bits),
    .io_data_1_out_valid(PE_605_io_data_1_out_valid),
    .io_data_1_out_bits(PE_605_io_data_1_out_bits),
    .io_data_0_in_valid(PE_605_io_data_0_in_valid),
    .io_data_0_in_bits(PE_605_io_data_0_in_bits),
    .io_data_0_out_valid(PE_605_io_data_0_out_valid),
    .io_data_0_out_bits(PE_605_io_data_0_out_bits)
  );
  PE PE_606 ( // @[pe.scala 187:13]
    .clock(PE_606_clock),
    .reset(PE_606_reset),
    .io_data_2_out_valid(PE_606_io_data_2_out_valid),
    .io_data_2_out_bits(PE_606_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_606_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_606_io_data_1_in_valid),
    .io_data_1_in_bits(PE_606_io_data_1_in_bits),
    .io_data_1_out_valid(PE_606_io_data_1_out_valid),
    .io_data_1_out_bits(PE_606_io_data_1_out_bits),
    .io_data_0_in_valid(PE_606_io_data_0_in_valid),
    .io_data_0_in_bits(PE_606_io_data_0_in_bits),
    .io_data_0_out_valid(PE_606_io_data_0_out_valid),
    .io_data_0_out_bits(PE_606_io_data_0_out_bits)
  );
  PE PE_607 ( // @[pe.scala 187:13]
    .clock(PE_607_clock),
    .reset(PE_607_reset),
    .io_data_2_out_valid(PE_607_io_data_2_out_valid),
    .io_data_2_out_bits(PE_607_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_607_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_607_io_data_1_in_valid),
    .io_data_1_in_bits(PE_607_io_data_1_in_bits),
    .io_data_1_out_valid(PE_607_io_data_1_out_valid),
    .io_data_1_out_bits(PE_607_io_data_1_out_bits),
    .io_data_0_in_valid(PE_607_io_data_0_in_valid),
    .io_data_0_in_bits(PE_607_io_data_0_in_bits),
    .io_data_0_out_valid(PE_607_io_data_0_out_valid),
    .io_data_0_out_bits(PE_607_io_data_0_out_bits)
  );
  PE PE_608 ( // @[pe.scala 187:13]
    .clock(PE_608_clock),
    .reset(PE_608_reset),
    .io_data_2_out_valid(PE_608_io_data_2_out_valid),
    .io_data_2_out_bits(PE_608_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_608_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_608_io_data_1_in_valid),
    .io_data_1_in_bits(PE_608_io_data_1_in_bits),
    .io_data_1_out_valid(PE_608_io_data_1_out_valid),
    .io_data_1_out_bits(PE_608_io_data_1_out_bits),
    .io_data_0_in_valid(PE_608_io_data_0_in_valid),
    .io_data_0_in_bits(PE_608_io_data_0_in_bits),
    .io_data_0_out_valid(PE_608_io_data_0_out_valid),
    .io_data_0_out_bits(PE_608_io_data_0_out_bits)
  );
  PE PE_609 ( // @[pe.scala 187:13]
    .clock(PE_609_clock),
    .reset(PE_609_reset),
    .io_data_2_out_valid(PE_609_io_data_2_out_valid),
    .io_data_2_out_bits(PE_609_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_609_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_609_io_data_1_in_valid),
    .io_data_1_in_bits(PE_609_io_data_1_in_bits),
    .io_data_1_out_valid(PE_609_io_data_1_out_valid),
    .io_data_1_out_bits(PE_609_io_data_1_out_bits),
    .io_data_0_in_valid(PE_609_io_data_0_in_valid),
    .io_data_0_in_bits(PE_609_io_data_0_in_bits),
    .io_data_0_out_valid(PE_609_io_data_0_out_valid),
    .io_data_0_out_bits(PE_609_io_data_0_out_bits)
  );
  PE PE_610 ( // @[pe.scala 187:13]
    .clock(PE_610_clock),
    .reset(PE_610_reset),
    .io_data_2_out_valid(PE_610_io_data_2_out_valid),
    .io_data_2_out_bits(PE_610_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_610_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_610_io_data_1_in_valid),
    .io_data_1_in_bits(PE_610_io_data_1_in_bits),
    .io_data_1_out_valid(PE_610_io_data_1_out_valid),
    .io_data_1_out_bits(PE_610_io_data_1_out_bits),
    .io_data_0_in_valid(PE_610_io_data_0_in_valid),
    .io_data_0_in_bits(PE_610_io_data_0_in_bits),
    .io_data_0_out_valid(PE_610_io_data_0_out_valid),
    .io_data_0_out_bits(PE_610_io_data_0_out_bits)
  );
  PE PE_611 ( // @[pe.scala 187:13]
    .clock(PE_611_clock),
    .reset(PE_611_reset),
    .io_data_2_out_valid(PE_611_io_data_2_out_valid),
    .io_data_2_out_bits(PE_611_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_611_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_611_io_data_1_in_valid),
    .io_data_1_in_bits(PE_611_io_data_1_in_bits),
    .io_data_1_out_valid(PE_611_io_data_1_out_valid),
    .io_data_1_out_bits(PE_611_io_data_1_out_bits),
    .io_data_0_in_valid(PE_611_io_data_0_in_valid),
    .io_data_0_in_bits(PE_611_io_data_0_in_bits),
    .io_data_0_out_valid(PE_611_io_data_0_out_valid),
    .io_data_0_out_bits(PE_611_io_data_0_out_bits)
  );
  PE PE_612 ( // @[pe.scala 187:13]
    .clock(PE_612_clock),
    .reset(PE_612_reset),
    .io_data_2_out_valid(PE_612_io_data_2_out_valid),
    .io_data_2_out_bits(PE_612_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_612_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_612_io_data_1_in_valid),
    .io_data_1_in_bits(PE_612_io_data_1_in_bits),
    .io_data_1_out_valid(PE_612_io_data_1_out_valid),
    .io_data_1_out_bits(PE_612_io_data_1_out_bits),
    .io_data_0_in_valid(PE_612_io_data_0_in_valid),
    .io_data_0_in_bits(PE_612_io_data_0_in_bits),
    .io_data_0_out_valid(PE_612_io_data_0_out_valid),
    .io_data_0_out_bits(PE_612_io_data_0_out_bits)
  );
  PE PE_613 ( // @[pe.scala 187:13]
    .clock(PE_613_clock),
    .reset(PE_613_reset),
    .io_data_2_out_valid(PE_613_io_data_2_out_valid),
    .io_data_2_out_bits(PE_613_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_613_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_613_io_data_1_in_valid),
    .io_data_1_in_bits(PE_613_io_data_1_in_bits),
    .io_data_1_out_valid(PE_613_io_data_1_out_valid),
    .io_data_1_out_bits(PE_613_io_data_1_out_bits),
    .io_data_0_in_valid(PE_613_io_data_0_in_valid),
    .io_data_0_in_bits(PE_613_io_data_0_in_bits),
    .io_data_0_out_valid(PE_613_io_data_0_out_valid),
    .io_data_0_out_bits(PE_613_io_data_0_out_bits)
  );
  PE PE_614 ( // @[pe.scala 187:13]
    .clock(PE_614_clock),
    .reset(PE_614_reset),
    .io_data_2_out_valid(PE_614_io_data_2_out_valid),
    .io_data_2_out_bits(PE_614_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_614_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_614_io_data_1_in_valid),
    .io_data_1_in_bits(PE_614_io_data_1_in_bits),
    .io_data_1_out_valid(PE_614_io_data_1_out_valid),
    .io_data_1_out_bits(PE_614_io_data_1_out_bits),
    .io_data_0_in_valid(PE_614_io_data_0_in_valid),
    .io_data_0_in_bits(PE_614_io_data_0_in_bits),
    .io_data_0_out_valid(PE_614_io_data_0_out_valid),
    .io_data_0_out_bits(PE_614_io_data_0_out_bits)
  );
  PE PE_615 ( // @[pe.scala 187:13]
    .clock(PE_615_clock),
    .reset(PE_615_reset),
    .io_data_2_out_valid(PE_615_io_data_2_out_valid),
    .io_data_2_out_bits(PE_615_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_615_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_615_io_data_1_in_valid),
    .io_data_1_in_bits(PE_615_io_data_1_in_bits),
    .io_data_1_out_valid(PE_615_io_data_1_out_valid),
    .io_data_1_out_bits(PE_615_io_data_1_out_bits),
    .io_data_0_in_valid(PE_615_io_data_0_in_valid),
    .io_data_0_in_bits(PE_615_io_data_0_in_bits),
    .io_data_0_out_valid(PE_615_io_data_0_out_valid),
    .io_data_0_out_bits(PE_615_io_data_0_out_bits)
  );
  PE PE_616 ( // @[pe.scala 187:13]
    .clock(PE_616_clock),
    .reset(PE_616_reset),
    .io_data_2_out_valid(PE_616_io_data_2_out_valid),
    .io_data_2_out_bits(PE_616_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_616_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_616_io_data_1_in_valid),
    .io_data_1_in_bits(PE_616_io_data_1_in_bits),
    .io_data_1_out_valid(PE_616_io_data_1_out_valid),
    .io_data_1_out_bits(PE_616_io_data_1_out_bits),
    .io_data_0_in_valid(PE_616_io_data_0_in_valid),
    .io_data_0_in_bits(PE_616_io_data_0_in_bits),
    .io_data_0_out_valid(PE_616_io_data_0_out_valid),
    .io_data_0_out_bits(PE_616_io_data_0_out_bits)
  );
  PE PE_617 ( // @[pe.scala 187:13]
    .clock(PE_617_clock),
    .reset(PE_617_reset),
    .io_data_2_out_valid(PE_617_io_data_2_out_valid),
    .io_data_2_out_bits(PE_617_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_617_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_617_io_data_1_in_valid),
    .io_data_1_in_bits(PE_617_io_data_1_in_bits),
    .io_data_1_out_valid(PE_617_io_data_1_out_valid),
    .io_data_1_out_bits(PE_617_io_data_1_out_bits),
    .io_data_0_in_valid(PE_617_io_data_0_in_valid),
    .io_data_0_in_bits(PE_617_io_data_0_in_bits),
    .io_data_0_out_valid(PE_617_io_data_0_out_valid),
    .io_data_0_out_bits(PE_617_io_data_0_out_bits)
  );
  PE PE_618 ( // @[pe.scala 187:13]
    .clock(PE_618_clock),
    .reset(PE_618_reset),
    .io_data_2_out_valid(PE_618_io_data_2_out_valid),
    .io_data_2_out_bits(PE_618_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_618_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_618_io_data_1_in_valid),
    .io_data_1_in_bits(PE_618_io_data_1_in_bits),
    .io_data_1_out_valid(PE_618_io_data_1_out_valid),
    .io_data_1_out_bits(PE_618_io_data_1_out_bits),
    .io_data_0_in_valid(PE_618_io_data_0_in_valid),
    .io_data_0_in_bits(PE_618_io_data_0_in_bits),
    .io_data_0_out_valid(PE_618_io_data_0_out_valid),
    .io_data_0_out_bits(PE_618_io_data_0_out_bits)
  );
  PE PE_619 ( // @[pe.scala 187:13]
    .clock(PE_619_clock),
    .reset(PE_619_reset),
    .io_data_2_out_valid(PE_619_io_data_2_out_valid),
    .io_data_2_out_bits(PE_619_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_619_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_619_io_data_1_in_valid),
    .io_data_1_in_bits(PE_619_io_data_1_in_bits),
    .io_data_1_out_valid(PE_619_io_data_1_out_valid),
    .io_data_1_out_bits(PE_619_io_data_1_out_bits),
    .io_data_0_in_valid(PE_619_io_data_0_in_valid),
    .io_data_0_in_bits(PE_619_io_data_0_in_bits),
    .io_data_0_out_valid(PE_619_io_data_0_out_valid),
    .io_data_0_out_bits(PE_619_io_data_0_out_bits)
  );
  PE PE_620 ( // @[pe.scala 187:13]
    .clock(PE_620_clock),
    .reset(PE_620_reset),
    .io_data_2_out_valid(PE_620_io_data_2_out_valid),
    .io_data_2_out_bits(PE_620_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_620_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_620_io_data_1_in_valid),
    .io_data_1_in_bits(PE_620_io_data_1_in_bits),
    .io_data_1_out_valid(PE_620_io_data_1_out_valid),
    .io_data_1_out_bits(PE_620_io_data_1_out_bits),
    .io_data_0_in_valid(PE_620_io_data_0_in_valid),
    .io_data_0_in_bits(PE_620_io_data_0_in_bits),
    .io_data_0_out_valid(PE_620_io_data_0_out_valid),
    .io_data_0_out_bits(PE_620_io_data_0_out_bits)
  );
  PE PE_621 ( // @[pe.scala 187:13]
    .clock(PE_621_clock),
    .reset(PE_621_reset),
    .io_data_2_out_valid(PE_621_io_data_2_out_valid),
    .io_data_2_out_bits(PE_621_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_621_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_621_io_data_1_in_valid),
    .io_data_1_in_bits(PE_621_io_data_1_in_bits),
    .io_data_1_out_valid(PE_621_io_data_1_out_valid),
    .io_data_1_out_bits(PE_621_io_data_1_out_bits),
    .io_data_0_in_valid(PE_621_io_data_0_in_valid),
    .io_data_0_in_bits(PE_621_io_data_0_in_bits),
    .io_data_0_out_valid(PE_621_io_data_0_out_valid),
    .io_data_0_out_bits(PE_621_io_data_0_out_bits)
  );
  PE PE_622 ( // @[pe.scala 187:13]
    .clock(PE_622_clock),
    .reset(PE_622_reset),
    .io_data_2_out_valid(PE_622_io_data_2_out_valid),
    .io_data_2_out_bits(PE_622_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_622_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_622_io_data_1_in_valid),
    .io_data_1_in_bits(PE_622_io_data_1_in_bits),
    .io_data_1_out_valid(PE_622_io_data_1_out_valid),
    .io_data_1_out_bits(PE_622_io_data_1_out_bits),
    .io_data_0_in_valid(PE_622_io_data_0_in_valid),
    .io_data_0_in_bits(PE_622_io_data_0_in_bits),
    .io_data_0_out_valid(PE_622_io_data_0_out_valid),
    .io_data_0_out_bits(PE_622_io_data_0_out_bits)
  );
  PE PE_623 ( // @[pe.scala 187:13]
    .clock(PE_623_clock),
    .reset(PE_623_reset),
    .io_data_2_out_valid(PE_623_io_data_2_out_valid),
    .io_data_2_out_bits(PE_623_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_623_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_623_io_data_1_in_valid),
    .io_data_1_in_bits(PE_623_io_data_1_in_bits),
    .io_data_1_out_valid(PE_623_io_data_1_out_valid),
    .io_data_1_out_bits(PE_623_io_data_1_out_bits),
    .io_data_0_in_valid(PE_623_io_data_0_in_valid),
    .io_data_0_in_bits(PE_623_io_data_0_in_bits),
    .io_data_0_out_valid(PE_623_io_data_0_out_valid),
    .io_data_0_out_bits(PE_623_io_data_0_out_bits)
  );
  PE PE_624 ( // @[pe.scala 187:13]
    .clock(PE_624_clock),
    .reset(PE_624_reset),
    .io_data_2_out_valid(PE_624_io_data_2_out_valid),
    .io_data_2_out_bits(PE_624_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_624_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_624_io_data_1_in_valid),
    .io_data_1_in_bits(PE_624_io_data_1_in_bits),
    .io_data_1_out_valid(PE_624_io_data_1_out_valid),
    .io_data_1_out_bits(PE_624_io_data_1_out_bits),
    .io_data_0_in_valid(PE_624_io_data_0_in_valid),
    .io_data_0_in_bits(PE_624_io_data_0_in_bits),
    .io_data_0_out_valid(PE_624_io_data_0_out_valid),
    .io_data_0_out_bits(PE_624_io_data_0_out_bits)
  );
  PE PE_625 ( // @[pe.scala 187:13]
    .clock(PE_625_clock),
    .reset(PE_625_reset),
    .io_data_2_out_valid(PE_625_io_data_2_out_valid),
    .io_data_2_out_bits(PE_625_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_625_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_625_io_data_1_in_valid),
    .io_data_1_in_bits(PE_625_io_data_1_in_bits),
    .io_data_1_out_valid(PE_625_io_data_1_out_valid),
    .io_data_1_out_bits(PE_625_io_data_1_out_bits),
    .io_data_0_in_valid(PE_625_io_data_0_in_valid),
    .io_data_0_in_bits(PE_625_io_data_0_in_bits),
    .io_data_0_out_valid(PE_625_io_data_0_out_valid),
    .io_data_0_out_bits(PE_625_io_data_0_out_bits)
  );
  PE PE_626 ( // @[pe.scala 187:13]
    .clock(PE_626_clock),
    .reset(PE_626_reset),
    .io_data_2_out_valid(PE_626_io_data_2_out_valid),
    .io_data_2_out_bits(PE_626_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_626_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_626_io_data_1_in_valid),
    .io_data_1_in_bits(PE_626_io_data_1_in_bits),
    .io_data_1_out_valid(PE_626_io_data_1_out_valid),
    .io_data_1_out_bits(PE_626_io_data_1_out_bits),
    .io_data_0_in_valid(PE_626_io_data_0_in_valid),
    .io_data_0_in_bits(PE_626_io_data_0_in_bits),
    .io_data_0_out_valid(PE_626_io_data_0_out_valid),
    .io_data_0_out_bits(PE_626_io_data_0_out_bits)
  );
  PE PE_627 ( // @[pe.scala 187:13]
    .clock(PE_627_clock),
    .reset(PE_627_reset),
    .io_data_2_out_valid(PE_627_io_data_2_out_valid),
    .io_data_2_out_bits(PE_627_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_627_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_627_io_data_1_in_valid),
    .io_data_1_in_bits(PE_627_io_data_1_in_bits),
    .io_data_1_out_valid(PE_627_io_data_1_out_valid),
    .io_data_1_out_bits(PE_627_io_data_1_out_bits),
    .io_data_0_in_valid(PE_627_io_data_0_in_valid),
    .io_data_0_in_bits(PE_627_io_data_0_in_bits),
    .io_data_0_out_valid(PE_627_io_data_0_out_valid),
    .io_data_0_out_bits(PE_627_io_data_0_out_bits)
  );
  PE PE_628 ( // @[pe.scala 187:13]
    .clock(PE_628_clock),
    .reset(PE_628_reset),
    .io_data_2_out_valid(PE_628_io_data_2_out_valid),
    .io_data_2_out_bits(PE_628_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_628_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_628_io_data_1_in_valid),
    .io_data_1_in_bits(PE_628_io_data_1_in_bits),
    .io_data_1_out_valid(PE_628_io_data_1_out_valid),
    .io_data_1_out_bits(PE_628_io_data_1_out_bits),
    .io_data_0_in_valid(PE_628_io_data_0_in_valid),
    .io_data_0_in_bits(PE_628_io_data_0_in_bits),
    .io_data_0_out_valid(PE_628_io_data_0_out_valid),
    .io_data_0_out_bits(PE_628_io_data_0_out_bits)
  );
  PE PE_629 ( // @[pe.scala 187:13]
    .clock(PE_629_clock),
    .reset(PE_629_reset),
    .io_data_2_out_valid(PE_629_io_data_2_out_valid),
    .io_data_2_out_bits(PE_629_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_629_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_629_io_data_1_in_valid),
    .io_data_1_in_bits(PE_629_io_data_1_in_bits),
    .io_data_1_out_valid(PE_629_io_data_1_out_valid),
    .io_data_1_out_bits(PE_629_io_data_1_out_bits),
    .io_data_0_in_valid(PE_629_io_data_0_in_valid),
    .io_data_0_in_bits(PE_629_io_data_0_in_bits),
    .io_data_0_out_valid(PE_629_io_data_0_out_valid),
    .io_data_0_out_bits(PE_629_io_data_0_out_bits)
  );
  PE PE_630 ( // @[pe.scala 187:13]
    .clock(PE_630_clock),
    .reset(PE_630_reset),
    .io_data_2_out_valid(PE_630_io_data_2_out_valid),
    .io_data_2_out_bits(PE_630_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_630_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_630_io_data_1_in_valid),
    .io_data_1_in_bits(PE_630_io_data_1_in_bits),
    .io_data_1_out_valid(PE_630_io_data_1_out_valid),
    .io_data_1_out_bits(PE_630_io_data_1_out_bits),
    .io_data_0_in_valid(PE_630_io_data_0_in_valid),
    .io_data_0_in_bits(PE_630_io_data_0_in_bits),
    .io_data_0_out_valid(PE_630_io_data_0_out_valid),
    .io_data_0_out_bits(PE_630_io_data_0_out_bits)
  );
  PE PE_631 ( // @[pe.scala 187:13]
    .clock(PE_631_clock),
    .reset(PE_631_reset),
    .io_data_2_out_valid(PE_631_io_data_2_out_valid),
    .io_data_2_out_bits(PE_631_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_631_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_631_io_data_1_in_valid),
    .io_data_1_in_bits(PE_631_io_data_1_in_bits),
    .io_data_1_out_valid(PE_631_io_data_1_out_valid),
    .io_data_1_out_bits(PE_631_io_data_1_out_bits),
    .io_data_0_in_valid(PE_631_io_data_0_in_valid),
    .io_data_0_in_bits(PE_631_io_data_0_in_bits),
    .io_data_0_out_valid(PE_631_io_data_0_out_valid),
    .io_data_0_out_bits(PE_631_io_data_0_out_bits)
  );
  PE PE_632 ( // @[pe.scala 187:13]
    .clock(PE_632_clock),
    .reset(PE_632_reset),
    .io_data_2_out_valid(PE_632_io_data_2_out_valid),
    .io_data_2_out_bits(PE_632_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_632_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_632_io_data_1_in_valid),
    .io_data_1_in_bits(PE_632_io_data_1_in_bits),
    .io_data_1_out_valid(PE_632_io_data_1_out_valid),
    .io_data_1_out_bits(PE_632_io_data_1_out_bits),
    .io_data_0_in_valid(PE_632_io_data_0_in_valid),
    .io_data_0_in_bits(PE_632_io_data_0_in_bits),
    .io_data_0_out_valid(PE_632_io_data_0_out_valid),
    .io_data_0_out_bits(PE_632_io_data_0_out_bits)
  );
  PE PE_633 ( // @[pe.scala 187:13]
    .clock(PE_633_clock),
    .reset(PE_633_reset),
    .io_data_2_out_valid(PE_633_io_data_2_out_valid),
    .io_data_2_out_bits(PE_633_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_633_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_633_io_data_1_in_valid),
    .io_data_1_in_bits(PE_633_io_data_1_in_bits),
    .io_data_1_out_valid(PE_633_io_data_1_out_valid),
    .io_data_1_out_bits(PE_633_io_data_1_out_bits),
    .io_data_0_in_valid(PE_633_io_data_0_in_valid),
    .io_data_0_in_bits(PE_633_io_data_0_in_bits),
    .io_data_0_out_valid(PE_633_io_data_0_out_valid),
    .io_data_0_out_bits(PE_633_io_data_0_out_bits)
  );
  PE PE_634 ( // @[pe.scala 187:13]
    .clock(PE_634_clock),
    .reset(PE_634_reset),
    .io_data_2_out_valid(PE_634_io_data_2_out_valid),
    .io_data_2_out_bits(PE_634_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_634_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_634_io_data_1_in_valid),
    .io_data_1_in_bits(PE_634_io_data_1_in_bits),
    .io_data_1_out_valid(PE_634_io_data_1_out_valid),
    .io_data_1_out_bits(PE_634_io_data_1_out_bits),
    .io_data_0_in_valid(PE_634_io_data_0_in_valid),
    .io_data_0_in_bits(PE_634_io_data_0_in_bits),
    .io_data_0_out_valid(PE_634_io_data_0_out_valid),
    .io_data_0_out_bits(PE_634_io_data_0_out_bits)
  );
  PE PE_635 ( // @[pe.scala 187:13]
    .clock(PE_635_clock),
    .reset(PE_635_reset),
    .io_data_2_out_valid(PE_635_io_data_2_out_valid),
    .io_data_2_out_bits(PE_635_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_635_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_635_io_data_1_in_valid),
    .io_data_1_in_bits(PE_635_io_data_1_in_bits),
    .io_data_1_out_valid(PE_635_io_data_1_out_valid),
    .io_data_1_out_bits(PE_635_io_data_1_out_bits),
    .io_data_0_in_valid(PE_635_io_data_0_in_valid),
    .io_data_0_in_bits(PE_635_io_data_0_in_bits),
    .io_data_0_out_valid(PE_635_io_data_0_out_valid),
    .io_data_0_out_bits(PE_635_io_data_0_out_bits)
  );
  PE PE_636 ( // @[pe.scala 187:13]
    .clock(PE_636_clock),
    .reset(PE_636_reset),
    .io_data_2_out_valid(PE_636_io_data_2_out_valid),
    .io_data_2_out_bits(PE_636_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_636_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_636_io_data_1_in_valid),
    .io_data_1_in_bits(PE_636_io_data_1_in_bits),
    .io_data_1_out_valid(PE_636_io_data_1_out_valid),
    .io_data_1_out_bits(PE_636_io_data_1_out_bits),
    .io_data_0_in_valid(PE_636_io_data_0_in_valid),
    .io_data_0_in_bits(PE_636_io_data_0_in_bits),
    .io_data_0_out_valid(PE_636_io_data_0_out_valid),
    .io_data_0_out_bits(PE_636_io_data_0_out_bits)
  );
  PE PE_637 ( // @[pe.scala 187:13]
    .clock(PE_637_clock),
    .reset(PE_637_reset),
    .io_data_2_out_valid(PE_637_io_data_2_out_valid),
    .io_data_2_out_bits(PE_637_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_637_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_637_io_data_1_in_valid),
    .io_data_1_in_bits(PE_637_io_data_1_in_bits),
    .io_data_1_out_valid(PE_637_io_data_1_out_valid),
    .io_data_1_out_bits(PE_637_io_data_1_out_bits),
    .io_data_0_in_valid(PE_637_io_data_0_in_valid),
    .io_data_0_in_bits(PE_637_io_data_0_in_bits),
    .io_data_0_out_valid(PE_637_io_data_0_out_valid),
    .io_data_0_out_bits(PE_637_io_data_0_out_bits)
  );
  PE PE_638 ( // @[pe.scala 187:13]
    .clock(PE_638_clock),
    .reset(PE_638_reset),
    .io_data_2_out_valid(PE_638_io_data_2_out_valid),
    .io_data_2_out_bits(PE_638_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_638_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_638_io_data_1_in_valid),
    .io_data_1_in_bits(PE_638_io_data_1_in_bits),
    .io_data_1_out_valid(PE_638_io_data_1_out_valid),
    .io_data_1_out_bits(PE_638_io_data_1_out_bits),
    .io_data_0_in_valid(PE_638_io_data_0_in_valid),
    .io_data_0_in_bits(PE_638_io_data_0_in_bits),
    .io_data_0_out_valid(PE_638_io_data_0_out_valid),
    .io_data_0_out_bits(PE_638_io_data_0_out_bits)
  );
  PE PE_639 ( // @[pe.scala 187:13]
    .clock(PE_639_clock),
    .reset(PE_639_reset),
    .io_data_2_out_valid(PE_639_io_data_2_out_valid),
    .io_data_2_out_bits(PE_639_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_639_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_639_io_data_1_in_valid),
    .io_data_1_in_bits(PE_639_io_data_1_in_bits),
    .io_data_1_out_valid(PE_639_io_data_1_out_valid),
    .io_data_1_out_bits(PE_639_io_data_1_out_bits),
    .io_data_0_in_valid(PE_639_io_data_0_in_valid),
    .io_data_0_in_bits(PE_639_io_data_0_in_bits),
    .io_data_0_out_valid(PE_639_io_data_0_out_valid),
    .io_data_0_out_bits(PE_639_io_data_0_out_bits)
  );
  PE PE_640 ( // @[pe.scala 187:13]
    .clock(PE_640_clock),
    .reset(PE_640_reset),
    .io_data_2_out_valid(PE_640_io_data_2_out_valid),
    .io_data_2_out_bits(PE_640_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_640_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_640_io_data_1_in_valid),
    .io_data_1_in_bits(PE_640_io_data_1_in_bits),
    .io_data_1_out_valid(PE_640_io_data_1_out_valid),
    .io_data_1_out_bits(PE_640_io_data_1_out_bits),
    .io_data_0_in_valid(PE_640_io_data_0_in_valid),
    .io_data_0_in_bits(PE_640_io_data_0_in_bits),
    .io_data_0_out_valid(PE_640_io_data_0_out_valid),
    .io_data_0_out_bits(PE_640_io_data_0_out_bits)
  );
  PE PE_641 ( // @[pe.scala 187:13]
    .clock(PE_641_clock),
    .reset(PE_641_reset),
    .io_data_2_out_valid(PE_641_io_data_2_out_valid),
    .io_data_2_out_bits(PE_641_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_641_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_641_io_data_1_in_valid),
    .io_data_1_in_bits(PE_641_io_data_1_in_bits),
    .io_data_1_out_valid(PE_641_io_data_1_out_valid),
    .io_data_1_out_bits(PE_641_io_data_1_out_bits),
    .io_data_0_in_valid(PE_641_io_data_0_in_valid),
    .io_data_0_in_bits(PE_641_io_data_0_in_bits),
    .io_data_0_out_valid(PE_641_io_data_0_out_valid),
    .io_data_0_out_bits(PE_641_io_data_0_out_bits)
  );
  PE PE_642 ( // @[pe.scala 187:13]
    .clock(PE_642_clock),
    .reset(PE_642_reset),
    .io_data_2_out_valid(PE_642_io_data_2_out_valid),
    .io_data_2_out_bits(PE_642_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_642_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_642_io_data_1_in_valid),
    .io_data_1_in_bits(PE_642_io_data_1_in_bits),
    .io_data_1_out_valid(PE_642_io_data_1_out_valid),
    .io_data_1_out_bits(PE_642_io_data_1_out_bits),
    .io_data_0_in_valid(PE_642_io_data_0_in_valid),
    .io_data_0_in_bits(PE_642_io_data_0_in_bits),
    .io_data_0_out_valid(PE_642_io_data_0_out_valid),
    .io_data_0_out_bits(PE_642_io_data_0_out_bits)
  );
  PE PE_643 ( // @[pe.scala 187:13]
    .clock(PE_643_clock),
    .reset(PE_643_reset),
    .io_data_2_out_valid(PE_643_io_data_2_out_valid),
    .io_data_2_out_bits(PE_643_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_643_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_643_io_data_1_in_valid),
    .io_data_1_in_bits(PE_643_io_data_1_in_bits),
    .io_data_1_out_valid(PE_643_io_data_1_out_valid),
    .io_data_1_out_bits(PE_643_io_data_1_out_bits),
    .io_data_0_in_valid(PE_643_io_data_0_in_valid),
    .io_data_0_in_bits(PE_643_io_data_0_in_bits),
    .io_data_0_out_valid(PE_643_io_data_0_out_valid),
    .io_data_0_out_bits(PE_643_io_data_0_out_bits)
  );
  PE PE_644 ( // @[pe.scala 187:13]
    .clock(PE_644_clock),
    .reset(PE_644_reset),
    .io_data_2_out_valid(PE_644_io_data_2_out_valid),
    .io_data_2_out_bits(PE_644_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_644_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_644_io_data_1_in_valid),
    .io_data_1_in_bits(PE_644_io_data_1_in_bits),
    .io_data_1_out_valid(PE_644_io_data_1_out_valid),
    .io_data_1_out_bits(PE_644_io_data_1_out_bits),
    .io_data_0_in_valid(PE_644_io_data_0_in_valid),
    .io_data_0_in_bits(PE_644_io_data_0_in_bits),
    .io_data_0_out_valid(PE_644_io_data_0_out_valid),
    .io_data_0_out_bits(PE_644_io_data_0_out_bits)
  );
  PE PE_645 ( // @[pe.scala 187:13]
    .clock(PE_645_clock),
    .reset(PE_645_reset),
    .io_data_2_out_valid(PE_645_io_data_2_out_valid),
    .io_data_2_out_bits(PE_645_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_645_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_645_io_data_1_in_valid),
    .io_data_1_in_bits(PE_645_io_data_1_in_bits),
    .io_data_1_out_valid(PE_645_io_data_1_out_valid),
    .io_data_1_out_bits(PE_645_io_data_1_out_bits),
    .io_data_0_in_valid(PE_645_io_data_0_in_valid),
    .io_data_0_in_bits(PE_645_io_data_0_in_bits),
    .io_data_0_out_valid(PE_645_io_data_0_out_valid),
    .io_data_0_out_bits(PE_645_io_data_0_out_bits)
  );
  PE PE_646 ( // @[pe.scala 187:13]
    .clock(PE_646_clock),
    .reset(PE_646_reset),
    .io_data_2_out_valid(PE_646_io_data_2_out_valid),
    .io_data_2_out_bits(PE_646_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_646_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_646_io_data_1_in_valid),
    .io_data_1_in_bits(PE_646_io_data_1_in_bits),
    .io_data_1_out_valid(PE_646_io_data_1_out_valid),
    .io_data_1_out_bits(PE_646_io_data_1_out_bits),
    .io_data_0_in_valid(PE_646_io_data_0_in_valid),
    .io_data_0_in_bits(PE_646_io_data_0_in_bits),
    .io_data_0_out_valid(PE_646_io_data_0_out_valid),
    .io_data_0_out_bits(PE_646_io_data_0_out_bits)
  );
  PE PE_647 ( // @[pe.scala 187:13]
    .clock(PE_647_clock),
    .reset(PE_647_reset),
    .io_data_2_out_valid(PE_647_io_data_2_out_valid),
    .io_data_2_out_bits(PE_647_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_647_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_647_io_data_1_in_valid),
    .io_data_1_in_bits(PE_647_io_data_1_in_bits),
    .io_data_1_out_valid(PE_647_io_data_1_out_valid),
    .io_data_1_out_bits(PE_647_io_data_1_out_bits),
    .io_data_0_in_valid(PE_647_io_data_0_in_valid),
    .io_data_0_in_bits(PE_647_io_data_0_in_bits),
    .io_data_0_out_valid(PE_647_io_data_0_out_valid),
    .io_data_0_out_bits(PE_647_io_data_0_out_bits)
  );
  PE PE_648 ( // @[pe.scala 187:13]
    .clock(PE_648_clock),
    .reset(PE_648_reset),
    .io_data_2_out_valid(PE_648_io_data_2_out_valid),
    .io_data_2_out_bits(PE_648_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_648_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_648_io_data_1_in_valid),
    .io_data_1_in_bits(PE_648_io_data_1_in_bits),
    .io_data_1_out_valid(PE_648_io_data_1_out_valid),
    .io_data_1_out_bits(PE_648_io_data_1_out_bits),
    .io_data_0_in_valid(PE_648_io_data_0_in_valid),
    .io_data_0_in_bits(PE_648_io_data_0_in_bits),
    .io_data_0_out_valid(PE_648_io_data_0_out_valid),
    .io_data_0_out_bits(PE_648_io_data_0_out_bits)
  );
  PE PE_649 ( // @[pe.scala 187:13]
    .clock(PE_649_clock),
    .reset(PE_649_reset),
    .io_data_2_out_valid(PE_649_io_data_2_out_valid),
    .io_data_2_out_bits(PE_649_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_649_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_649_io_data_1_in_valid),
    .io_data_1_in_bits(PE_649_io_data_1_in_bits),
    .io_data_1_out_valid(PE_649_io_data_1_out_valid),
    .io_data_1_out_bits(PE_649_io_data_1_out_bits),
    .io_data_0_in_valid(PE_649_io_data_0_in_valid),
    .io_data_0_in_bits(PE_649_io_data_0_in_bits),
    .io_data_0_out_valid(PE_649_io_data_0_out_valid),
    .io_data_0_out_bits(PE_649_io_data_0_out_bits)
  );
  PE PE_650 ( // @[pe.scala 187:13]
    .clock(PE_650_clock),
    .reset(PE_650_reset),
    .io_data_2_out_valid(PE_650_io_data_2_out_valid),
    .io_data_2_out_bits(PE_650_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_650_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_650_io_data_1_in_valid),
    .io_data_1_in_bits(PE_650_io_data_1_in_bits),
    .io_data_1_out_valid(PE_650_io_data_1_out_valid),
    .io_data_1_out_bits(PE_650_io_data_1_out_bits),
    .io_data_0_in_valid(PE_650_io_data_0_in_valid),
    .io_data_0_in_bits(PE_650_io_data_0_in_bits),
    .io_data_0_out_valid(PE_650_io_data_0_out_valid),
    .io_data_0_out_bits(PE_650_io_data_0_out_bits)
  );
  PE PE_651 ( // @[pe.scala 187:13]
    .clock(PE_651_clock),
    .reset(PE_651_reset),
    .io_data_2_out_valid(PE_651_io_data_2_out_valid),
    .io_data_2_out_bits(PE_651_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_651_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_651_io_data_1_in_valid),
    .io_data_1_in_bits(PE_651_io_data_1_in_bits),
    .io_data_1_out_valid(PE_651_io_data_1_out_valid),
    .io_data_1_out_bits(PE_651_io_data_1_out_bits),
    .io_data_0_in_valid(PE_651_io_data_0_in_valid),
    .io_data_0_in_bits(PE_651_io_data_0_in_bits),
    .io_data_0_out_valid(PE_651_io_data_0_out_valid),
    .io_data_0_out_bits(PE_651_io_data_0_out_bits)
  );
  PE PE_652 ( // @[pe.scala 187:13]
    .clock(PE_652_clock),
    .reset(PE_652_reset),
    .io_data_2_out_valid(PE_652_io_data_2_out_valid),
    .io_data_2_out_bits(PE_652_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_652_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_652_io_data_1_in_valid),
    .io_data_1_in_bits(PE_652_io_data_1_in_bits),
    .io_data_1_out_valid(PE_652_io_data_1_out_valid),
    .io_data_1_out_bits(PE_652_io_data_1_out_bits),
    .io_data_0_in_valid(PE_652_io_data_0_in_valid),
    .io_data_0_in_bits(PE_652_io_data_0_in_bits),
    .io_data_0_out_valid(PE_652_io_data_0_out_valid),
    .io_data_0_out_bits(PE_652_io_data_0_out_bits)
  );
  PE PE_653 ( // @[pe.scala 187:13]
    .clock(PE_653_clock),
    .reset(PE_653_reset),
    .io_data_2_out_valid(PE_653_io_data_2_out_valid),
    .io_data_2_out_bits(PE_653_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_653_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_653_io_data_1_in_valid),
    .io_data_1_in_bits(PE_653_io_data_1_in_bits),
    .io_data_1_out_valid(PE_653_io_data_1_out_valid),
    .io_data_1_out_bits(PE_653_io_data_1_out_bits),
    .io_data_0_in_valid(PE_653_io_data_0_in_valid),
    .io_data_0_in_bits(PE_653_io_data_0_in_bits),
    .io_data_0_out_valid(PE_653_io_data_0_out_valid),
    .io_data_0_out_bits(PE_653_io_data_0_out_bits)
  );
  PE PE_654 ( // @[pe.scala 187:13]
    .clock(PE_654_clock),
    .reset(PE_654_reset),
    .io_data_2_out_valid(PE_654_io_data_2_out_valid),
    .io_data_2_out_bits(PE_654_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_654_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_654_io_data_1_in_valid),
    .io_data_1_in_bits(PE_654_io_data_1_in_bits),
    .io_data_1_out_valid(PE_654_io_data_1_out_valid),
    .io_data_1_out_bits(PE_654_io_data_1_out_bits),
    .io_data_0_in_valid(PE_654_io_data_0_in_valid),
    .io_data_0_in_bits(PE_654_io_data_0_in_bits),
    .io_data_0_out_valid(PE_654_io_data_0_out_valid),
    .io_data_0_out_bits(PE_654_io_data_0_out_bits)
  );
  PE PE_655 ( // @[pe.scala 187:13]
    .clock(PE_655_clock),
    .reset(PE_655_reset),
    .io_data_2_out_valid(PE_655_io_data_2_out_valid),
    .io_data_2_out_bits(PE_655_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_655_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_655_io_data_1_in_valid),
    .io_data_1_in_bits(PE_655_io_data_1_in_bits),
    .io_data_1_out_valid(PE_655_io_data_1_out_valid),
    .io_data_1_out_bits(PE_655_io_data_1_out_bits),
    .io_data_0_in_valid(PE_655_io_data_0_in_valid),
    .io_data_0_in_bits(PE_655_io_data_0_in_bits),
    .io_data_0_out_valid(PE_655_io_data_0_out_valid),
    .io_data_0_out_bits(PE_655_io_data_0_out_bits)
  );
  PE PE_656 ( // @[pe.scala 187:13]
    .clock(PE_656_clock),
    .reset(PE_656_reset),
    .io_data_2_out_valid(PE_656_io_data_2_out_valid),
    .io_data_2_out_bits(PE_656_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_656_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_656_io_data_1_in_valid),
    .io_data_1_in_bits(PE_656_io_data_1_in_bits),
    .io_data_1_out_valid(PE_656_io_data_1_out_valid),
    .io_data_1_out_bits(PE_656_io_data_1_out_bits),
    .io_data_0_in_valid(PE_656_io_data_0_in_valid),
    .io_data_0_in_bits(PE_656_io_data_0_in_bits),
    .io_data_0_out_valid(PE_656_io_data_0_out_valid),
    .io_data_0_out_bits(PE_656_io_data_0_out_bits)
  );
  PE PE_657 ( // @[pe.scala 187:13]
    .clock(PE_657_clock),
    .reset(PE_657_reset),
    .io_data_2_out_valid(PE_657_io_data_2_out_valid),
    .io_data_2_out_bits(PE_657_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_657_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_657_io_data_1_in_valid),
    .io_data_1_in_bits(PE_657_io_data_1_in_bits),
    .io_data_1_out_valid(PE_657_io_data_1_out_valid),
    .io_data_1_out_bits(PE_657_io_data_1_out_bits),
    .io_data_0_in_valid(PE_657_io_data_0_in_valid),
    .io_data_0_in_bits(PE_657_io_data_0_in_bits),
    .io_data_0_out_valid(PE_657_io_data_0_out_valid),
    .io_data_0_out_bits(PE_657_io_data_0_out_bits)
  );
  PE PE_658 ( // @[pe.scala 187:13]
    .clock(PE_658_clock),
    .reset(PE_658_reset),
    .io_data_2_out_valid(PE_658_io_data_2_out_valid),
    .io_data_2_out_bits(PE_658_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_658_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_658_io_data_1_in_valid),
    .io_data_1_in_bits(PE_658_io_data_1_in_bits),
    .io_data_1_out_valid(PE_658_io_data_1_out_valid),
    .io_data_1_out_bits(PE_658_io_data_1_out_bits),
    .io_data_0_in_valid(PE_658_io_data_0_in_valid),
    .io_data_0_in_bits(PE_658_io_data_0_in_bits),
    .io_data_0_out_valid(PE_658_io_data_0_out_valid),
    .io_data_0_out_bits(PE_658_io_data_0_out_bits)
  );
  PE PE_659 ( // @[pe.scala 187:13]
    .clock(PE_659_clock),
    .reset(PE_659_reset),
    .io_data_2_out_valid(PE_659_io_data_2_out_valid),
    .io_data_2_out_bits(PE_659_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_659_io_data_2_sig_stat2trans),
    .io_data_1_in_valid(PE_659_io_data_1_in_valid),
    .io_data_1_in_bits(PE_659_io_data_1_in_bits),
    .io_data_1_out_valid(PE_659_io_data_1_out_valid),
    .io_data_1_out_bits(PE_659_io_data_1_out_bits),
    .io_data_0_in_valid(PE_659_io_data_0_in_valid),
    .io_data_0_in_bits(PE_659_io_data_0_in_bits),
    .io_data_0_out_valid(PE_659_io_data_0_out_valid),
    .io_data_0_out_bits(PE_659_io_data_0_out_bits)
  );
  PENetwork PENetwork ( // @[pe.scala 229:13]
    .io_to_pes_0_in_valid(PENetwork_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_io_to_pes_15_out_bits),
    .io_to_pes_16_in_valid(PENetwork_io_to_pes_16_in_valid),
    .io_to_pes_16_in_bits(PENetwork_io_to_pes_16_in_bits),
    .io_to_pes_16_out_valid(PENetwork_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_io_to_pes_16_out_bits),
    .io_to_pes_17_in_valid(PENetwork_io_to_pes_17_in_valid),
    .io_to_pes_17_in_bits(PENetwork_io_to_pes_17_in_bits),
    .io_to_pes_17_out_valid(PENetwork_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_io_to_pes_17_out_bits),
    .io_to_pes_18_in_valid(PENetwork_io_to_pes_18_in_valid),
    .io_to_pes_18_in_bits(PENetwork_io_to_pes_18_in_bits),
    .io_to_pes_18_out_valid(PENetwork_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_io_to_pes_18_out_bits),
    .io_to_pes_19_in_valid(PENetwork_io_to_pes_19_in_valid),
    .io_to_pes_19_in_bits(PENetwork_io_to_pes_19_in_bits),
    .io_to_pes_19_out_valid(PENetwork_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_io_to_pes_19_out_bits),
    .io_to_pes_20_in_valid(PENetwork_io_to_pes_20_in_valid),
    .io_to_pes_20_in_bits(PENetwork_io_to_pes_20_in_bits),
    .io_to_pes_20_out_valid(PENetwork_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_io_to_pes_20_out_bits),
    .io_to_pes_21_in_valid(PENetwork_io_to_pes_21_in_valid),
    .io_to_pes_21_in_bits(PENetwork_io_to_pes_21_in_bits),
    .io_to_pes_21_out_valid(PENetwork_io_to_pes_21_out_valid),
    .io_to_pes_21_out_bits(PENetwork_io_to_pes_21_out_bits),
    .io_to_pes_22_in_valid(PENetwork_io_to_pes_22_in_valid),
    .io_to_pes_22_in_bits(PENetwork_io_to_pes_22_in_bits),
    .io_to_pes_22_out_valid(PENetwork_io_to_pes_22_out_valid),
    .io_to_pes_22_out_bits(PENetwork_io_to_pes_22_out_bits),
    .io_to_pes_23_in_valid(PENetwork_io_to_pes_23_in_valid),
    .io_to_pes_23_in_bits(PENetwork_io_to_pes_23_in_bits),
    .io_to_pes_23_out_valid(PENetwork_io_to_pes_23_out_valid),
    .io_to_pes_23_out_bits(PENetwork_io_to_pes_23_out_bits),
    .io_to_pes_24_in_valid(PENetwork_io_to_pes_24_in_valid),
    .io_to_pes_24_in_bits(PENetwork_io_to_pes_24_in_bits),
    .io_to_pes_24_out_valid(PENetwork_io_to_pes_24_out_valid),
    .io_to_pes_24_out_bits(PENetwork_io_to_pes_24_out_bits),
    .io_to_pes_25_in_valid(PENetwork_io_to_pes_25_in_valid),
    .io_to_pes_25_in_bits(PENetwork_io_to_pes_25_in_bits),
    .io_to_pes_25_out_valid(PENetwork_io_to_pes_25_out_valid),
    .io_to_pes_25_out_bits(PENetwork_io_to_pes_25_out_bits),
    .io_to_pes_26_in_valid(PENetwork_io_to_pes_26_in_valid),
    .io_to_pes_26_in_bits(PENetwork_io_to_pes_26_in_bits),
    .io_to_pes_26_out_valid(PENetwork_io_to_pes_26_out_valid),
    .io_to_pes_26_out_bits(PENetwork_io_to_pes_26_out_bits),
    .io_to_pes_27_in_valid(PENetwork_io_to_pes_27_in_valid),
    .io_to_pes_27_in_bits(PENetwork_io_to_pes_27_in_bits),
    .io_to_pes_27_out_valid(PENetwork_io_to_pes_27_out_valid),
    .io_to_pes_27_out_bits(PENetwork_io_to_pes_27_out_bits),
    .io_to_pes_28_in_valid(PENetwork_io_to_pes_28_in_valid),
    .io_to_pes_28_in_bits(PENetwork_io_to_pes_28_in_bits),
    .io_to_pes_28_out_valid(PENetwork_io_to_pes_28_out_valid),
    .io_to_pes_28_out_bits(PENetwork_io_to_pes_28_out_bits),
    .io_to_pes_29_in_valid(PENetwork_io_to_pes_29_in_valid),
    .io_to_pes_29_in_bits(PENetwork_io_to_pes_29_in_bits),
    .io_to_mem_valid(PENetwork_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_io_to_mem_bits)
  );
  PENetwork PENetwork_1 ( // @[pe.scala 229:13]
    .io_to_pes_0_in_valid(PENetwork_1_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_1_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_1_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_1_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_1_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_1_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_1_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_1_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_1_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_1_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_1_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_1_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_1_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_1_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_1_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_1_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_1_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_1_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_1_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_1_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_1_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_1_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_1_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_1_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_1_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_1_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_1_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_1_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_1_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_1_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_1_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_1_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_1_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_1_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_1_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_1_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_1_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_1_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_1_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_1_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_1_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_1_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_1_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_1_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_1_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_1_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_1_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_1_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_1_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_1_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_1_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_1_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_1_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_1_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_1_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_1_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_1_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_1_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_1_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_1_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_1_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_1_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_1_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_1_io_to_pes_15_out_bits),
    .io_to_pes_16_in_valid(PENetwork_1_io_to_pes_16_in_valid),
    .io_to_pes_16_in_bits(PENetwork_1_io_to_pes_16_in_bits),
    .io_to_pes_16_out_valid(PENetwork_1_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_1_io_to_pes_16_out_bits),
    .io_to_pes_17_in_valid(PENetwork_1_io_to_pes_17_in_valid),
    .io_to_pes_17_in_bits(PENetwork_1_io_to_pes_17_in_bits),
    .io_to_pes_17_out_valid(PENetwork_1_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_1_io_to_pes_17_out_bits),
    .io_to_pes_18_in_valid(PENetwork_1_io_to_pes_18_in_valid),
    .io_to_pes_18_in_bits(PENetwork_1_io_to_pes_18_in_bits),
    .io_to_pes_18_out_valid(PENetwork_1_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_1_io_to_pes_18_out_bits),
    .io_to_pes_19_in_valid(PENetwork_1_io_to_pes_19_in_valid),
    .io_to_pes_19_in_bits(PENetwork_1_io_to_pes_19_in_bits),
    .io_to_pes_19_out_valid(PENetwork_1_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_1_io_to_pes_19_out_bits),
    .io_to_pes_20_in_valid(PENetwork_1_io_to_pes_20_in_valid),
    .io_to_pes_20_in_bits(PENetwork_1_io_to_pes_20_in_bits),
    .io_to_pes_20_out_valid(PENetwork_1_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_1_io_to_pes_20_out_bits),
    .io_to_pes_21_in_valid(PENetwork_1_io_to_pes_21_in_valid),
    .io_to_pes_21_in_bits(PENetwork_1_io_to_pes_21_in_bits),
    .io_to_pes_21_out_valid(PENetwork_1_io_to_pes_21_out_valid),
    .io_to_pes_21_out_bits(PENetwork_1_io_to_pes_21_out_bits),
    .io_to_pes_22_in_valid(PENetwork_1_io_to_pes_22_in_valid),
    .io_to_pes_22_in_bits(PENetwork_1_io_to_pes_22_in_bits),
    .io_to_pes_22_out_valid(PENetwork_1_io_to_pes_22_out_valid),
    .io_to_pes_22_out_bits(PENetwork_1_io_to_pes_22_out_bits),
    .io_to_pes_23_in_valid(PENetwork_1_io_to_pes_23_in_valid),
    .io_to_pes_23_in_bits(PENetwork_1_io_to_pes_23_in_bits),
    .io_to_pes_23_out_valid(PENetwork_1_io_to_pes_23_out_valid),
    .io_to_pes_23_out_bits(PENetwork_1_io_to_pes_23_out_bits),
    .io_to_pes_24_in_valid(PENetwork_1_io_to_pes_24_in_valid),
    .io_to_pes_24_in_bits(PENetwork_1_io_to_pes_24_in_bits),
    .io_to_pes_24_out_valid(PENetwork_1_io_to_pes_24_out_valid),
    .io_to_pes_24_out_bits(PENetwork_1_io_to_pes_24_out_bits),
    .io_to_pes_25_in_valid(PENetwork_1_io_to_pes_25_in_valid),
    .io_to_pes_25_in_bits(PENetwork_1_io_to_pes_25_in_bits),
    .io_to_pes_25_out_valid(PENetwork_1_io_to_pes_25_out_valid),
    .io_to_pes_25_out_bits(PENetwork_1_io_to_pes_25_out_bits),
    .io_to_pes_26_in_valid(PENetwork_1_io_to_pes_26_in_valid),
    .io_to_pes_26_in_bits(PENetwork_1_io_to_pes_26_in_bits),
    .io_to_pes_26_out_valid(PENetwork_1_io_to_pes_26_out_valid),
    .io_to_pes_26_out_bits(PENetwork_1_io_to_pes_26_out_bits),
    .io_to_pes_27_in_valid(PENetwork_1_io_to_pes_27_in_valid),
    .io_to_pes_27_in_bits(PENetwork_1_io_to_pes_27_in_bits),
    .io_to_pes_27_out_valid(PENetwork_1_io_to_pes_27_out_valid),
    .io_to_pes_27_out_bits(PENetwork_1_io_to_pes_27_out_bits),
    .io_to_pes_28_in_valid(PENetwork_1_io_to_pes_28_in_valid),
    .io_to_pes_28_in_bits(PENetwork_1_io_to_pes_28_in_bits),
    .io_to_pes_28_out_valid(PENetwork_1_io_to_pes_28_out_valid),
    .io_to_pes_28_out_bits(PENetwork_1_io_to_pes_28_out_bits),
    .io_to_pes_29_in_valid(PENetwork_1_io_to_pes_29_in_valid),
    .io_to_pes_29_in_bits(PENetwork_1_io_to_pes_29_in_bits),
    .io_to_mem_valid(PENetwork_1_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_1_io_to_mem_bits)
  );
  PENetwork PENetwork_2 ( // @[pe.scala 229:13]
    .io_to_pes_0_in_valid(PENetwork_2_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_2_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_2_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_2_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_2_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_2_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_2_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_2_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_2_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_2_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_2_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_2_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_2_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_2_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_2_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_2_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_2_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_2_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_2_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_2_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_2_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_2_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_2_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_2_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_2_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_2_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_2_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_2_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_2_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_2_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_2_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_2_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_2_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_2_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_2_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_2_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_2_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_2_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_2_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_2_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_2_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_2_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_2_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_2_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_2_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_2_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_2_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_2_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_2_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_2_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_2_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_2_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_2_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_2_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_2_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_2_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_2_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_2_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_2_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_2_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_2_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_2_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_2_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_2_io_to_pes_15_out_bits),
    .io_to_pes_16_in_valid(PENetwork_2_io_to_pes_16_in_valid),
    .io_to_pes_16_in_bits(PENetwork_2_io_to_pes_16_in_bits),
    .io_to_pes_16_out_valid(PENetwork_2_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_2_io_to_pes_16_out_bits),
    .io_to_pes_17_in_valid(PENetwork_2_io_to_pes_17_in_valid),
    .io_to_pes_17_in_bits(PENetwork_2_io_to_pes_17_in_bits),
    .io_to_pes_17_out_valid(PENetwork_2_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_2_io_to_pes_17_out_bits),
    .io_to_pes_18_in_valid(PENetwork_2_io_to_pes_18_in_valid),
    .io_to_pes_18_in_bits(PENetwork_2_io_to_pes_18_in_bits),
    .io_to_pes_18_out_valid(PENetwork_2_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_2_io_to_pes_18_out_bits),
    .io_to_pes_19_in_valid(PENetwork_2_io_to_pes_19_in_valid),
    .io_to_pes_19_in_bits(PENetwork_2_io_to_pes_19_in_bits),
    .io_to_pes_19_out_valid(PENetwork_2_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_2_io_to_pes_19_out_bits),
    .io_to_pes_20_in_valid(PENetwork_2_io_to_pes_20_in_valid),
    .io_to_pes_20_in_bits(PENetwork_2_io_to_pes_20_in_bits),
    .io_to_pes_20_out_valid(PENetwork_2_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_2_io_to_pes_20_out_bits),
    .io_to_pes_21_in_valid(PENetwork_2_io_to_pes_21_in_valid),
    .io_to_pes_21_in_bits(PENetwork_2_io_to_pes_21_in_bits),
    .io_to_pes_21_out_valid(PENetwork_2_io_to_pes_21_out_valid),
    .io_to_pes_21_out_bits(PENetwork_2_io_to_pes_21_out_bits),
    .io_to_pes_22_in_valid(PENetwork_2_io_to_pes_22_in_valid),
    .io_to_pes_22_in_bits(PENetwork_2_io_to_pes_22_in_bits),
    .io_to_pes_22_out_valid(PENetwork_2_io_to_pes_22_out_valid),
    .io_to_pes_22_out_bits(PENetwork_2_io_to_pes_22_out_bits),
    .io_to_pes_23_in_valid(PENetwork_2_io_to_pes_23_in_valid),
    .io_to_pes_23_in_bits(PENetwork_2_io_to_pes_23_in_bits),
    .io_to_pes_23_out_valid(PENetwork_2_io_to_pes_23_out_valid),
    .io_to_pes_23_out_bits(PENetwork_2_io_to_pes_23_out_bits),
    .io_to_pes_24_in_valid(PENetwork_2_io_to_pes_24_in_valid),
    .io_to_pes_24_in_bits(PENetwork_2_io_to_pes_24_in_bits),
    .io_to_pes_24_out_valid(PENetwork_2_io_to_pes_24_out_valid),
    .io_to_pes_24_out_bits(PENetwork_2_io_to_pes_24_out_bits),
    .io_to_pes_25_in_valid(PENetwork_2_io_to_pes_25_in_valid),
    .io_to_pes_25_in_bits(PENetwork_2_io_to_pes_25_in_bits),
    .io_to_pes_25_out_valid(PENetwork_2_io_to_pes_25_out_valid),
    .io_to_pes_25_out_bits(PENetwork_2_io_to_pes_25_out_bits),
    .io_to_pes_26_in_valid(PENetwork_2_io_to_pes_26_in_valid),
    .io_to_pes_26_in_bits(PENetwork_2_io_to_pes_26_in_bits),
    .io_to_pes_26_out_valid(PENetwork_2_io_to_pes_26_out_valid),
    .io_to_pes_26_out_bits(PENetwork_2_io_to_pes_26_out_bits),
    .io_to_pes_27_in_valid(PENetwork_2_io_to_pes_27_in_valid),
    .io_to_pes_27_in_bits(PENetwork_2_io_to_pes_27_in_bits),
    .io_to_pes_27_out_valid(PENetwork_2_io_to_pes_27_out_valid),
    .io_to_pes_27_out_bits(PENetwork_2_io_to_pes_27_out_bits),
    .io_to_pes_28_in_valid(PENetwork_2_io_to_pes_28_in_valid),
    .io_to_pes_28_in_bits(PENetwork_2_io_to_pes_28_in_bits),
    .io_to_pes_28_out_valid(PENetwork_2_io_to_pes_28_out_valid),
    .io_to_pes_28_out_bits(PENetwork_2_io_to_pes_28_out_bits),
    .io_to_pes_29_in_valid(PENetwork_2_io_to_pes_29_in_valid),
    .io_to_pes_29_in_bits(PENetwork_2_io_to_pes_29_in_bits),
    .io_to_mem_valid(PENetwork_2_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_2_io_to_mem_bits)
  );
  PENetwork PENetwork_3 ( // @[pe.scala 229:13]
    .io_to_pes_0_in_valid(PENetwork_3_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_3_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_3_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_3_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_3_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_3_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_3_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_3_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_3_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_3_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_3_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_3_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_3_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_3_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_3_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_3_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_3_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_3_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_3_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_3_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_3_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_3_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_3_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_3_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_3_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_3_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_3_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_3_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_3_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_3_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_3_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_3_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_3_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_3_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_3_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_3_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_3_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_3_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_3_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_3_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_3_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_3_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_3_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_3_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_3_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_3_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_3_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_3_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_3_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_3_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_3_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_3_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_3_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_3_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_3_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_3_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_3_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_3_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_3_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_3_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_3_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_3_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_3_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_3_io_to_pes_15_out_bits),
    .io_to_pes_16_in_valid(PENetwork_3_io_to_pes_16_in_valid),
    .io_to_pes_16_in_bits(PENetwork_3_io_to_pes_16_in_bits),
    .io_to_pes_16_out_valid(PENetwork_3_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_3_io_to_pes_16_out_bits),
    .io_to_pes_17_in_valid(PENetwork_3_io_to_pes_17_in_valid),
    .io_to_pes_17_in_bits(PENetwork_3_io_to_pes_17_in_bits),
    .io_to_pes_17_out_valid(PENetwork_3_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_3_io_to_pes_17_out_bits),
    .io_to_pes_18_in_valid(PENetwork_3_io_to_pes_18_in_valid),
    .io_to_pes_18_in_bits(PENetwork_3_io_to_pes_18_in_bits),
    .io_to_pes_18_out_valid(PENetwork_3_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_3_io_to_pes_18_out_bits),
    .io_to_pes_19_in_valid(PENetwork_3_io_to_pes_19_in_valid),
    .io_to_pes_19_in_bits(PENetwork_3_io_to_pes_19_in_bits),
    .io_to_pes_19_out_valid(PENetwork_3_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_3_io_to_pes_19_out_bits),
    .io_to_pes_20_in_valid(PENetwork_3_io_to_pes_20_in_valid),
    .io_to_pes_20_in_bits(PENetwork_3_io_to_pes_20_in_bits),
    .io_to_pes_20_out_valid(PENetwork_3_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_3_io_to_pes_20_out_bits),
    .io_to_pes_21_in_valid(PENetwork_3_io_to_pes_21_in_valid),
    .io_to_pes_21_in_bits(PENetwork_3_io_to_pes_21_in_bits),
    .io_to_pes_21_out_valid(PENetwork_3_io_to_pes_21_out_valid),
    .io_to_pes_21_out_bits(PENetwork_3_io_to_pes_21_out_bits),
    .io_to_pes_22_in_valid(PENetwork_3_io_to_pes_22_in_valid),
    .io_to_pes_22_in_bits(PENetwork_3_io_to_pes_22_in_bits),
    .io_to_pes_22_out_valid(PENetwork_3_io_to_pes_22_out_valid),
    .io_to_pes_22_out_bits(PENetwork_3_io_to_pes_22_out_bits),
    .io_to_pes_23_in_valid(PENetwork_3_io_to_pes_23_in_valid),
    .io_to_pes_23_in_bits(PENetwork_3_io_to_pes_23_in_bits),
    .io_to_pes_23_out_valid(PENetwork_3_io_to_pes_23_out_valid),
    .io_to_pes_23_out_bits(PENetwork_3_io_to_pes_23_out_bits),
    .io_to_pes_24_in_valid(PENetwork_3_io_to_pes_24_in_valid),
    .io_to_pes_24_in_bits(PENetwork_3_io_to_pes_24_in_bits),
    .io_to_pes_24_out_valid(PENetwork_3_io_to_pes_24_out_valid),
    .io_to_pes_24_out_bits(PENetwork_3_io_to_pes_24_out_bits),
    .io_to_pes_25_in_valid(PENetwork_3_io_to_pes_25_in_valid),
    .io_to_pes_25_in_bits(PENetwork_3_io_to_pes_25_in_bits),
    .io_to_pes_25_out_valid(PENetwork_3_io_to_pes_25_out_valid),
    .io_to_pes_25_out_bits(PENetwork_3_io_to_pes_25_out_bits),
    .io_to_pes_26_in_valid(PENetwork_3_io_to_pes_26_in_valid),
    .io_to_pes_26_in_bits(PENetwork_3_io_to_pes_26_in_bits),
    .io_to_pes_26_out_valid(PENetwork_3_io_to_pes_26_out_valid),
    .io_to_pes_26_out_bits(PENetwork_3_io_to_pes_26_out_bits),
    .io_to_pes_27_in_valid(PENetwork_3_io_to_pes_27_in_valid),
    .io_to_pes_27_in_bits(PENetwork_3_io_to_pes_27_in_bits),
    .io_to_pes_27_out_valid(PENetwork_3_io_to_pes_27_out_valid),
    .io_to_pes_27_out_bits(PENetwork_3_io_to_pes_27_out_bits),
    .io_to_pes_28_in_valid(PENetwork_3_io_to_pes_28_in_valid),
    .io_to_pes_28_in_bits(PENetwork_3_io_to_pes_28_in_bits),
    .io_to_pes_28_out_valid(PENetwork_3_io_to_pes_28_out_valid),
    .io_to_pes_28_out_bits(PENetwork_3_io_to_pes_28_out_bits),
    .io_to_pes_29_in_valid(PENetwork_3_io_to_pes_29_in_valid),
    .io_to_pes_29_in_bits(PENetwork_3_io_to_pes_29_in_bits),
    .io_to_mem_valid(PENetwork_3_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_3_io_to_mem_bits)
  );
  PENetwork PENetwork_4 ( // @[pe.scala 229:13]
    .io_to_pes_0_in_valid(PENetwork_4_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_4_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_4_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_4_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_4_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_4_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_4_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_4_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_4_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_4_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_4_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_4_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_4_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_4_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_4_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_4_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_4_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_4_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_4_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_4_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_4_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_4_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_4_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_4_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_4_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_4_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_4_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_4_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_4_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_4_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_4_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_4_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_4_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_4_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_4_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_4_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_4_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_4_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_4_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_4_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_4_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_4_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_4_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_4_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_4_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_4_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_4_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_4_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_4_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_4_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_4_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_4_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_4_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_4_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_4_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_4_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_4_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_4_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_4_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_4_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_4_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_4_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_4_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_4_io_to_pes_15_out_bits),
    .io_to_pes_16_in_valid(PENetwork_4_io_to_pes_16_in_valid),
    .io_to_pes_16_in_bits(PENetwork_4_io_to_pes_16_in_bits),
    .io_to_pes_16_out_valid(PENetwork_4_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_4_io_to_pes_16_out_bits),
    .io_to_pes_17_in_valid(PENetwork_4_io_to_pes_17_in_valid),
    .io_to_pes_17_in_bits(PENetwork_4_io_to_pes_17_in_bits),
    .io_to_pes_17_out_valid(PENetwork_4_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_4_io_to_pes_17_out_bits),
    .io_to_pes_18_in_valid(PENetwork_4_io_to_pes_18_in_valid),
    .io_to_pes_18_in_bits(PENetwork_4_io_to_pes_18_in_bits),
    .io_to_pes_18_out_valid(PENetwork_4_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_4_io_to_pes_18_out_bits),
    .io_to_pes_19_in_valid(PENetwork_4_io_to_pes_19_in_valid),
    .io_to_pes_19_in_bits(PENetwork_4_io_to_pes_19_in_bits),
    .io_to_pes_19_out_valid(PENetwork_4_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_4_io_to_pes_19_out_bits),
    .io_to_pes_20_in_valid(PENetwork_4_io_to_pes_20_in_valid),
    .io_to_pes_20_in_bits(PENetwork_4_io_to_pes_20_in_bits),
    .io_to_pes_20_out_valid(PENetwork_4_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_4_io_to_pes_20_out_bits),
    .io_to_pes_21_in_valid(PENetwork_4_io_to_pes_21_in_valid),
    .io_to_pes_21_in_bits(PENetwork_4_io_to_pes_21_in_bits),
    .io_to_pes_21_out_valid(PENetwork_4_io_to_pes_21_out_valid),
    .io_to_pes_21_out_bits(PENetwork_4_io_to_pes_21_out_bits),
    .io_to_pes_22_in_valid(PENetwork_4_io_to_pes_22_in_valid),
    .io_to_pes_22_in_bits(PENetwork_4_io_to_pes_22_in_bits),
    .io_to_pes_22_out_valid(PENetwork_4_io_to_pes_22_out_valid),
    .io_to_pes_22_out_bits(PENetwork_4_io_to_pes_22_out_bits),
    .io_to_pes_23_in_valid(PENetwork_4_io_to_pes_23_in_valid),
    .io_to_pes_23_in_bits(PENetwork_4_io_to_pes_23_in_bits),
    .io_to_pes_23_out_valid(PENetwork_4_io_to_pes_23_out_valid),
    .io_to_pes_23_out_bits(PENetwork_4_io_to_pes_23_out_bits),
    .io_to_pes_24_in_valid(PENetwork_4_io_to_pes_24_in_valid),
    .io_to_pes_24_in_bits(PENetwork_4_io_to_pes_24_in_bits),
    .io_to_pes_24_out_valid(PENetwork_4_io_to_pes_24_out_valid),
    .io_to_pes_24_out_bits(PENetwork_4_io_to_pes_24_out_bits),
    .io_to_pes_25_in_valid(PENetwork_4_io_to_pes_25_in_valid),
    .io_to_pes_25_in_bits(PENetwork_4_io_to_pes_25_in_bits),
    .io_to_pes_25_out_valid(PENetwork_4_io_to_pes_25_out_valid),
    .io_to_pes_25_out_bits(PENetwork_4_io_to_pes_25_out_bits),
    .io_to_pes_26_in_valid(PENetwork_4_io_to_pes_26_in_valid),
    .io_to_pes_26_in_bits(PENetwork_4_io_to_pes_26_in_bits),
    .io_to_pes_26_out_valid(PENetwork_4_io_to_pes_26_out_valid),
    .io_to_pes_26_out_bits(PENetwork_4_io_to_pes_26_out_bits),
    .io_to_pes_27_in_valid(PENetwork_4_io_to_pes_27_in_valid),
    .io_to_pes_27_in_bits(PENetwork_4_io_to_pes_27_in_bits),
    .io_to_pes_27_out_valid(PENetwork_4_io_to_pes_27_out_valid),
    .io_to_pes_27_out_bits(PENetwork_4_io_to_pes_27_out_bits),
    .io_to_pes_28_in_valid(PENetwork_4_io_to_pes_28_in_valid),
    .io_to_pes_28_in_bits(PENetwork_4_io_to_pes_28_in_bits),
    .io_to_pes_28_out_valid(PENetwork_4_io_to_pes_28_out_valid),
    .io_to_pes_28_out_bits(PENetwork_4_io_to_pes_28_out_bits),
    .io_to_pes_29_in_valid(PENetwork_4_io_to_pes_29_in_valid),
    .io_to_pes_29_in_bits(PENetwork_4_io_to_pes_29_in_bits),
    .io_to_mem_valid(PENetwork_4_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_4_io_to_mem_bits)
  );
  PENetwork PENetwork_5 ( // @[pe.scala 229:13]
    .io_to_pes_0_in_valid(PENetwork_5_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_5_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_5_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_5_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_5_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_5_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_5_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_5_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_5_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_5_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_5_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_5_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_5_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_5_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_5_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_5_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_5_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_5_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_5_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_5_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_5_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_5_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_5_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_5_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_5_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_5_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_5_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_5_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_5_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_5_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_5_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_5_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_5_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_5_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_5_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_5_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_5_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_5_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_5_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_5_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_5_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_5_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_5_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_5_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_5_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_5_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_5_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_5_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_5_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_5_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_5_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_5_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_5_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_5_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_5_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_5_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_5_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_5_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_5_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_5_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_5_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_5_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_5_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_5_io_to_pes_15_out_bits),
    .io_to_pes_16_in_valid(PENetwork_5_io_to_pes_16_in_valid),
    .io_to_pes_16_in_bits(PENetwork_5_io_to_pes_16_in_bits),
    .io_to_pes_16_out_valid(PENetwork_5_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_5_io_to_pes_16_out_bits),
    .io_to_pes_17_in_valid(PENetwork_5_io_to_pes_17_in_valid),
    .io_to_pes_17_in_bits(PENetwork_5_io_to_pes_17_in_bits),
    .io_to_pes_17_out_valid(PENetwork_5_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_5_io_to_pes_17_out_bits),
    .io_to_pes_18_in_valid(PENetwork_5_io_to_pes_18_in_valid),
    .io_to_pes_18_in_bits(PENetwork_5_io_to_pes_18_in_bits),
    .io_to_pes_18_out_valid(PENetwork_5_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_5_io_to_pes_18_out_bits),
    .io_to_pes_19_in_valid(PENetwork_5_io_to_pes_19_in_valid),
    .io_to_pes_19_in_bits(PENetwork_5_io_to_pes_19_in_bits),
    .io_to_pes_19_out_valid(PENetwork_5_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_5_io_to_pes_19_out_bits),
    .io_to_pes_20_in_valid(PENetwork_5_io_to_pes_20_in_valid),
    .io_to_pes_20_in_bits(PENetwork_5_io_to_pes_20_in_bits),
    .io_to_pes_20_out_valid(PENetwork_5_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_5_io_to_pes_20_out_bits),
    .io_to_pes_21_in_valid(PENetwork_5_io_to_pes_21_in_valid),
    .io_to_pes_21_in_bits(PENetwork_5_io_to_pes_21_in_bits),
    .io_to_pes_21_out_valid(PENetwork_5_io_to_pes_21_out_valid),
    .io_to_pes_21_out_bits(PENetwork_5_io_to_pes_21_out_bits),
    .io_to_pes_22_in_valid(PENetwork_5_io_to_pes_22_in_valid),
    .io_to_pes_22_in_bits(PENetwork_5_io_to_pes_22_in_bits),
    .io_to_pes_22_out_valid(PENetwork_5_io_to_pes_22_out_valid),
    .io_to_pes_22_out_bits(PENetwork_5_io_to_pes_22_out_bits),
    .io_to_pes_23_in_valid(PENetwork_5_io_to_pes_23_in_valid),
    .io_to_pes_23_in_bits(PENetwork_5_io_to_pes_23_in_bits),
    .io_to_pes_23_out_valid(PENetwork_5_io_to_pes_23_out_valid),
    .io_to_pes_23_out_bits(PENetwork_5_io_to_pes_23_out_bits),
    .io_to_pes_24_in_valid(PENetwork_5_io_to_pes_24_in_valid),
    .io_to_pes_24_in_bits(PENetwork_5_io_to_pes_24_in_bits),
    .io_to_pes_24_out_valid(PENetwork_5_io_to_pes_24_out_valid),
    .io_to_pes_24_out_bits(PENetwork_5_io_to_pes_24_out_bits),
    .io_to_pes_25_in_valid(PENetwork_5_io_to_pes_25_in_valid),
    .io_to_pes_25_in_bits(PENetwork_5_io_to_pes_25_in_bits),
    .io_to_pes_25_out_valid(PENetwork_5_io_to_pes_25_out_valid),
    .io_to_pes_25_out_bits(PENetwork_5_io_to_pes_25_out_bits),
    .io_to_pes_26_in_valid(PENetwork_5_io_to_pes_26_in_valid),
    .io_to_pes_26_in_bits(PENetwork_5_io_to_pes_26_in_bits),
    .io_to_pes_26_out_valid(PENetwork_5_io_to_pes_26_out_valid),
    .io_to_pes_26_out_bits(PENetwork_5_io_to_pes_26_out_bits),
    .io_to_pes_27_in_valid(PENetwork_5_io_to_pes_27_in_valid),
    .io_to_pes_27_in_bits(PENetwork_5_io_to_pes_27_in_bits),
    .io_to_pes_27_out_valid(PENetwork_5_io_to_pes_27_out_valid),
    .io_to_pes_27_out_bits(PENetwork_5_io_to_pes_27_out_bits),
    .io_to_pes_28_in_valid(PENetwork_5_io_to_pes_28_in_valid),
    .io_to_pes_28_in_bits(PENetwork_5_io_to_pes_28_in_bits),
    .io_to_pes_28_out_valid(PENetwork_5_io_to_pes_28_out_valid),
    .io_to_pes_28_out_bits(PENetwork_5_io_to_pes_28_out_bits),
    .io_to_pes_29_in_valid(PENetwork_5_io_to_pes_29_in_valid),
    .io_to_pes_29_in_bits(PENetwork_5_io_to_pes_29_in_bits),
    .io_to_mem_valid(PENetwork_5_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_5_io_to_mem_bits)
  );
  PENetwork PENetwork_6 ( // @[pe.scala 229:13]
    .io_to_pes_0_in_valid(PENetwork_6_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_6_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_6_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_6_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_6_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_6_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_6_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_6_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_6_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_6_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_6_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_6_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_6_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_6_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_6_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_6_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_6_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_6_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_6_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_6_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_6_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_6_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_6_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_6_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_6_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_6_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_6_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_6_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_6_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_6_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_6_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_6_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_6_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_6_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_6_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_6_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_6_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_6_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_6_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_6_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_6_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_6_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_6_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_6_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_6_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_6_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_6_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_6_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_6_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_6_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_6_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_6_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_6_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_6_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_6_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_6_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_6_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_6_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_6_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_6_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_6_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_6_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_6_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_6_io_to_pes_15_out_bits),
    .io_to_pes_16_in_valid(PENetwork_6_io_to_pes_16_in_valid),
    .io_to_pes_16_in_bits(PENetwork_6_io_to_pes_16_in_bits),
    .io_to_pes_16_out_valid(PENetwork_6_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_6_io_to_pes_16_out_bits),
    .io_to_pes_17_in_valid(PENetwork_6_io_to_pes_17_in_valid),
    .io_to_pes_17_in_bits(PENetwork_6_io_to_pes_17_in_bits),
    .io_to_pes_17_out_valid(PENetwork_6_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_6_io_to_pes_17_out_bits),
    .io_to_pes_18_in_valid(PENetwork_6_io_to_pes_18_in_valid),
    .io_to_pes_18_in_bits(PENetwork_6_io_to_pes_18_in_bits),
    .io_to_pes_18_out_valid(PENetwork_6_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_6_io_to_pes_18_out_bits),
    .io_to_pes_19_in_valid(PENetwork_6_io_to_pes_19_in_valid),
    .io_to_pes_19_in_bits(PENetwork_6_io_to_pes_19_in_bits),
    .io_to_pes_19_out_valid(PENetwork_6_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_6_io_to_pes_19_out_bits),
    .io_to_pes_20_in_valid(PENetwork_6_io_to_pes_20_in_valid),
    .io_to_pes_20_in_bits(PENetwork_6_io_to_pes_20_in_bits),
    .io_to_pes_20_out_valid(PENetwork_6_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_6_io_to_pes_20_out_bits),
    .io_to_pes_21_in_valid(PENetwork_6_io_to_pes_21_in_valid),
    .io_to_pes_21_in_bits(PENetwork_6_io_to_pes_21_in_bits),
    .io_to_pes_21_out_valid(PENetwork_6_io_to_pes_21_out_valid),
    .io_to_pes_21_out_bits(PENetwork_6_io_to_pes_21_out_bits),
    .io_to_pes_22_in_valid(PENetwork_6_io_to_pes_22_in_valid),
    .io_to_pes_22_in_bits(PENetwork_6_io_to_pes_22_in_bits),
    .io_to_pes_22_out_valid(PENetwork_6_io_to_pes_22_out_valid),
    .io_to_pes_22_out_bits(PENetwork_6_io_to_pes_22_out_bits),
    .io_to_pes_23_in_valid(PENetwork_6_io_to_pes_23_in_valid),
    .io_to_pes_23_in_bits(PENetwork_6_io_to_pes_23_in_bits),
    .io_to_pes_23_out_valid(PENetwork_6_io_to_pes_23_out_valid),
    .io_to_pes_23_out_bits(PENetwork_6_io_to_pes_23_out_bits),
    .io_to_pes_24_in_valid(PENetwork_6_io_to_pes_24_in_valid),
    .io_to_pes_24_in_bits(PENetwork_6_io_to_pes_24_in_bits),
    .io_to_pes_24_out_valid(PENetwork_6_io_to_pes_24_out_valid),
    .io_to_pes_24_out_bits(PENetwork_6_io_to_pes_24_out_bits),
    .io_to_pes_25_in_valid(PENetwork_6_io_to_pes_25_in_valid),
    .io_to_pes_25_in_bits(PENetwork_6_io_to_pes_25_in_bits),
    .io_to_pes_25_out_valid(PENetwork_6_io_to_pes_25_out_valid),
    .io_to_pes_25_out_bits(PENetwork_6_io_to_pes_25_out_bits),
    .io_to_pes_26_in_valid(PENetwork_6_io_to_pes_26_in_valid),
    .io_to_pes_26_in_bits(PENetwork_6_io_to_pes_26_in_bits),
    .io_to_pes_26_out_valid(PENetwork_6_io_to_pes_26_out_valid),
    .io_to_pes_26_out_bits(PENetwork_6_io_to_pes_26_out_bits),
    .io_to_pes_27_in_valid(PENetwork_6_io_to_pes_27_in_valid),
    .io_to_pes_27_in_bits(PENetwork_6_io_to_pes_27_in_bits),
    .io_to_pes_27_out_valid(PENetwork_6_io_to_pes_27_out_valid),
    .io_to_pes_27_out_bits(PENetwork_6_io_to_pes_27_out_bits),
    .io_to_pes_28_in_valid(PENetwork_6_io_to_pes_28_in_valid),
    .io_to_pes_28_in_bits(PENetwork_6_io_to_pes_28_in_bits),
    .io_to_pes_28_out_valid(PENetwork_6_io_to_pes_28_out_valid),
    .io_to_pes_28_out_bits(PENetwork_6_io_to_pes_28_out_bits),
    .io_to_pes_29_in_valid(PENetwork_6_io_to_pes_29_in_valid),
    .io_to_pes_29_in_bits(PENetwork_6_io_to_pes_29_in_bits),
    .io_to_mem_valid(PENetwork_6_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_6_io_to_mem_bits)
  );
  PENetwork PENetwork_7 ( // @[pe.scala 229:13]
    .io_to_pes_0_in_valid(PENetwork_7_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_7_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_7_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_7_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_7_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_7_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_7_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_7_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_7_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_7_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_7_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_7_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_7_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_7_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_7_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_7_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_7_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_7_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_7_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_7_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_7_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_7_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_7_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_7_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_7_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_7_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_7_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_7_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_7_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_7_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_7_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_7_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_7_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_7_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_7_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_7_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_7_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_7_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_7_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_7_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_7_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_7_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_7_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_7_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_7_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_7_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_7_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_7_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_7_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_7_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_7_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_7_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_7_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_7_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_7_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_7_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_7_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_7_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_7_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_7_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_7_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_7_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_7_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_7_io_to_pes_15_out_bits),
    .io_to_pes_16_in_valid(PENetwork_7_io_to_pes_16_in_valid),
    .io_to_pes_16_in_bits(PENetwork_7_io_to_pes_16_in_bits),
    .io_to_pes_16_out_valid(PENetwork_7_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_7_io_to_pes_16_out_bits),
    .io_to_pes_17_in_valid(PENetwork_7_io_to_pes_17_in_valid),
    .io_to_pes_17_in_bits(PENetwork_7_io_to_pes_17_in_bits),
    .io_to_pes_17_out_valid(PENetwork_7_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_7_io_to_pes_17_out_bits),
    .io_to_pes_18_in_valid(PENetwork_7_io_to_pes_18_in_valid),
    .io_to_pes_18_in_bits(PENetwork_7_io_to_pes_18_in_bits),
    .io_to_pes_18_out_valid(PENetwork_7_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_7_io_to_pes_18_out_bits),
    .io_to_pes_19_in_valid(PENetwork_7_io_to_pes_19_in_valid),
    .io_to_pes_19_in_bits(PENetwork_7_io_to_pes_19_in_bits),
    .io_to_pes_19_out_valid(PENetwork_7_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_7_io_to_pes_19_out_bits),
    .io_to_pes_20_in_valid(PENetwork_7_io_to_pes_20_in_valid),
    .io_to_pes_20_in_bits(PENetwork_7_io_to_pes_20_in_bits),
    .io_to_pes_20_out_valid(PENetwork_7_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_7_io_to_pes_20_out_bits),
    .io_to_pes_21_in_valid(PENetwork_7_io_to_pes_21_in_valid),
    .io_to_pes_21_in_bits(PENetwork_7_io_to_pes_21_in_bits),
    .io_to_pes_21_out_valid(PENetwork_7_io_to_pes_21_out_valid),
    .io_to_pes_21_out_bits(PENetwork_7_io_to_pes_21_out_bits),
    .io_to_pes_22_in_valid(PENetwork_7_io_to_pes_22_in_valid),
    .io_to_pes_22_in_bits(PENetwork_7_io_to_pes_22_in_bits),
    .io_to_pes_22_out_valid(PENetwork_7_io_to_pes_22_out_valid),
    .io_to_pes_22_out_bits(PENetwork_7_io_to_pes_22_out_bits),
    .io_to_pes_23_in_valid(PENetwork_7_io_to_pes_23_in_valid),
    .io_to_pes_23_in_bits(PENetwork_7_io_to_pes_23_in_bits),
    .io_to_pes_23_out_valid(PENetwork_7_io_to_pes_23_out_valid),
    .io_to_pes_23_out_bits(PENetwork_7_io_to_pes_23_out_bits),
    .io_to_pes_24_in_valid(PENetwork_7_io_to_pes_24_in_valid),
    .io_to_pes_24_in_bits(PENetwork_7_io_to_pes_24_in_bits),
    .io_to_pes_24_out_valid(PENetwork_7_io_to_pes_24_out_valid),
    .io_to_pes_24_out_bits(PENetwork_7_io_to_pes_24_out_bits),
    .io_to_pes_25_in_valid(PENetwork_7_io_to_pes_25_in_valid),
    .io_to_pes_25_in_bits(PENetwork_7_io_to_pes_25_in_bits),
    .io_to_pes_25_out_valid(PENetwork_7_io_to_pes_25_out_valid),
    .io_to_pes_25_out_bits(PENetwork_7_io_to_pes_25_out_bits),
    .io_to_pes_26_in_valid(PENetwork_7_io_to_pes_26_in_valid),
    .io_to_pes_26_in_bits(PENetwork_7_io_to_pes_26_in_bits),
    .io_to_pes_26_out_valid(PENetwork_7_io_to_pes_26_out_valid),
    .io_to_pes_26_out_bits(PENetwork_7_io_to_pes_26_out_bits),
    .io_to_pes_27_in_valid(PENetwork_7_io_to_pes_27_in_valid),
    .io_to_pes_27_in_bits(PENetwork_7_io_to_pes_27_in_bits),
    .io_to_pes_27_out_valid(PENetwork_7_io_to_pes_27_out_valid),
    .io_to_pes_27_out_bits(PENetwork_7_io_to_pes_27_out_bits),
    .io_to_pes_28_in_valid(PENetwork_7_io_to_pes_28_in_valid),
    .io_to_pes_28_in_bits(PENetwork_7_io_to_pes_28_in_bits),
    .io_to_pes_28_out_valid(PENetwork_7_io_to_pes_28_out_valid),
    .io_to_pes_28_out_bits(PENetwork_7_io_to_pes_28_out_bits),
    .io_to_pes_29_in_valid(PENetwork_7_io_to_pes_29_in_valid),
    .io_to_pes_29_in_bits(PENetwork_7_io_to_pes_29_in_bits),
    .io_to_mem_valid(PENetwork_7_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_7_io_to_mem_bits)
  );
  PENetwork PENetwork_8 ( // @[pe.scala 229:13]
    .io_to_pes_0_in_valid(PENetwork_8_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_8_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_8_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_8_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_8_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_8_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_8_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_8_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_8_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_8_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_8_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_8_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_8_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_8_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_8_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_8_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_8_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_8_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_8_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_8_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_8_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_8_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_8_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_8_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_8_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_8_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_8_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_8_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_8_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_8_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_8_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_8_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_8_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_8_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_8_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_8_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_8_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_8_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_8_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_8_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_8_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_8_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_8_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_8_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_8_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_8_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_8_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_8_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_8_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_8_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_8_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_8_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_8_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_8_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_8_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_8_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_8_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_8_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_8_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_8_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_8_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_8_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_8_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_8_io_to_pes_15_out_bits),
    .io_to_pes_16_in_valid(PENetwork_8_io_to_pes_16_in_valid),
    .io_to_pes_16_in_bits(PENetwork_8_io_to_pes_16_in_bits),
    .io_to_pes_16_out_valid(PENetwork_8_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_8_io_to_pes_16_out_bits),
    .io_to_pes_17_in_valid(PENetwork_8_io_to_pes_17_in_valid),
    .io_to_pes_17_in_bits(PENetwork_8_io_to_pes_17_in_bits),
    .io_to_pes_17_out_valid(PENetwork_8_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_8_io_to_pes_17_out_bits),
    .io_to_pes_18_in_valid(PENetwork_8_io_to_pes_18_in_valid),
    .io_to_pes_18_in_bits(PENetwork_8_io_to_pes_18_in_bits),
    .io_to_pes_18_out_valid(PENetwork_8_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_8_io_to_pes_18_out_bits),
    .io_to_pes_19_in_valid(PENetwork_8_io_to_pes_19_in_valid),
    .io_to_pes_19_in_bits(PENetwork_8_io_to_pes_19_in_bits),
    .io_to_pes_19_out_valid(PENetwork_8_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_8_io_to_pes_19_out_bits),
    .io_to_pes_20_in_valid(PENetwork_8_io_to_pes_20_in_valid),
    .io_to_pes_20_in_bits(PENetwork_8_io_to_pes_20_in_bits),
    .io_to_pes_20_out_valid(PENetwork_8_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_8_io_to_pes_20_out_bits),
    .io_to_pes_21_in_valid(PENetwork_8_io_to_pes_21_in_valid),
    .io_to_pes_21_in_bits(PENetwork_8_io_to_pes_21_in_bits),
    .io_to_pes_21_out_valid(PENetwork_8_io_to_pes_21_out_valid),
    .io_to_pes_21_out_bits(PENetwork_8_io_to_pes_21_out_bits),
    .io_to_pes_22_in_valid(PENetwork_8_io_to_pes_22_in_valid),
    .io_to_pes_22_in_bits(PENetwork_8_io_to_pes_22_in_bits),
    .io_to_pes_22_out_valid(PENetwork_8_io_to_pes_22_out_valid),
    .io_to_pes_22_out_bits(PENetwork_8_io_to_pes_22_out_bits),
    .io_to_pes_23_in_valid(PENetwork_8_io_to_pes_23_in_valid),
    .io_to_pes_23_in_bits(PENetwork_8_io_to_pes_23_in_bits),
    .io_to_pes_23_out_valid(PENetwork_8_io_to_pes_23_out_valid),
    .io_to_pes_23_out_bits(PENetwork_8_io_to_pes_23_out_bits),
    .io_to_pes_24_in_valid(PENetwork_8_io_to_pes_24_in_valid),
    .io_to_pes_24_in_bits(PENetwork_8_io_to_pes_24_in_bits),
    .io_to_pes_24_out_valid(PENetwork_8_io_to_pes_24_out_valid),
    .io_to_pes_24_out_bits(PENetwork_8_io_to_pes_24_out_bits),
    .io_to_pes_25_in_valid(PENetwork_8_io_to_pes_25_in_valid),
    .io_to_pes_25_in_bits(PENetwork_8_io_to_pes_25_in_bits),
    .io_to_pes_25_out_valid(PENetwork_8_io_to_pes_25_out_valid),
    .io_to_pes_25_out_bits(PENetwork_8_io_to_pes_25_out_bits),
    .io_to_pes_26_in_valid(PENetwork_8_io_to_pes_26_in_valid),
    .io_to_pes_26_in_bits(PENetwork_8_io_to_pes_26_in_bits),
    .io_to_pes_26_out_valid(PENetwork_8_io_to_pes_26_out_valid),
    .io_to_pes_26_out_bits(PENetwork_8_io_to_pes_26_out_bits),
    .io_to_pes_27_in_valid(PENetwork_8_io_to_pes_27_in_valid),
    .io_to_pes_27_in_bits(PENetwork_8_io_to_pes_27_in_bits),
    .io_to_pes_27_out_valid(PENetwork_8_io_to_pes_27_out_valid),
    .io_to_pes_27_out_bits(PENetwork_8_io_to_pes_27_out_bits),
    .io_to_pes_28_in_valid(PENetwork_8_io_to_pes_28_in_valid),
    .io_to_pes_28_in_bits(PENetwork_8_io_to_pes_28_in_bits),
    .io_to_pes_28_out_valid(PENetwork_8_io_to_pes_28_out_valid),
    .io_to_pes_28_out_bits(PENetwork_8_io_to_pes_28_out_bits),
    .io_to_pes_29_in_valid(PENetwork_8_io_to_pes_29_in_valid),
    .io_to_pes_29_in_bits(PENetwork_8_io_to_pes_29_in_bits),
    .io_to_mem_valid(PENetwork_8_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_8_io_to_mem_bits)
  );
  PENetwork PENetwork_9 ( // @[pe.scala 229:13]
    .io_to_pes_0_in_valid(PENetwork_9_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_9_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_9_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_9_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_9_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_9_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_9_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_9_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_9_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_9_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_9_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_9_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_9_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_9_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_9_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_9_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_9_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_9_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_9_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_9_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_9_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_9_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_9_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_9_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_9_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_9_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_9_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_9_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_9_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_9_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_9_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_9_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_9_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_9_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_9_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_9_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_9_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_9_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_9_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_9_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_9_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_9_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_9_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_9_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_9_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_9_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_9_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_9_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_9_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_9_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_9_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_9_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_9_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_9_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_9_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_9_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_9_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_9_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_9_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_9_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_9_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_9_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_9_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_9_io_to_pes_15_out_bits),
    .io_to_pes_16_in_valid(PENetwork_9_io_to_pes_16_in_valid),
    .io_to_pes_16_in_bits(PENetwork_9_io_to_pes_16_in_bits),
    .io_to_pes_16_out_valid(PENetwork_9_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_9_io_to_pes_16_out_bits),
    .io_to_pes_17_in_valid(PENetwork_9_io_to_pes_17_in_valid),
    .io_to_pes_17_in_bits(PENetwork_9_io_to_pes_17_in_bits),
    .io_to_pes_17_out_valid(PENetwork_9_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_9_io_to_pes_17_out_bits),
    .io_to_pes_18_in_valid(PENetwork_9_io_to_pes_18_in_valid),
    .io_to_pes_18_in_bits(PENetwork_9_io_to_pes_18_in_bits),
    .io_to_pes_18_out_valid(PENetwork_9_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_9_io_to_pes_18_out_bits),
    .io_to_pes_19_in_valid(PENetwork_9_io_to_pes_19_in_valid),
    .io_to_pes_19_in_bits(PENetwork_9_io_to_pes_19_in_bits),
    .io_to_pes_19_out_valid(PENetwork_9_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_9_io_to_pes_19_out_bits),
    .io_to_pes_20_in_valid(PENetwork_9_io_to_pes_20_in_valid),
    .io_to_pes_20_in_bits(PENetwork_9_io_to_pes_20_in_bits),
    .io_to_pes_20_out_valid(PENetwork_9_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_9_io_to_pes_20_out_bits),
    .io_to_pes_21_in_valid(PENetwork_9_io_to_pes_21_in_valid),
    .io_to_pes_21_in_bits(PENetwork_9_io_to_pes_21_in_bits),
    .io_to_pes_21_out_valid(PENetwork_9_io_to_pes_21_out_valid),
    .io_to_pes_21_out_bits(PENetwork_9_io_to_pes_21_out_bits),
    .io_to_pes_22_in_valid(PENetwork_9_io_to_pes_22_in_valid),
    .io_to_pes_22_in_bits(PENetwork_9_io_to_pes_22_in_bits),
    .io_to_pes_22_out_valid(PENetwork_9_io_to_pes_22_out_valid),
    .io_to_pes_22_out_bits(PENetwork_9_io_to_pes_22_out_bits),
    .io_to_pes_23_in_valid(PENetwork_9_io_to_pes_23_in_valid),
    .io_to_pes_23_in_bits(PENetwork_9_io_to_pes_23_in_bits),
    .io_to_pes_23_out_valid(PENetwork_9_io_to_pes_23_out_valid),
    .io_to_pes_23_out_bits(PENetwork_9_io_to_pes_23_out_bits),
    .io_to_pes_24_in_valid(PENetwork_9_io_to_pes_24_in_valid),
    .io_to_pes_24_in_bits(PENetwork_9_io_to_pes_24_in_bits),
    .io_to_pes_24_out_valid(PENetwork_9_io_to_pes_24_out_valid),
    .io_to_pes_24_out_bits(PENetwork_9_io_to_pes_24_out_bits),
    .io_to_pes_25_in_valid(PENetwork_9_io_to_pes_25_in_valid),
    .io_to_pes_25_in_bits(PENetwork_9_io_to_pes_25_in_bits),
    .io_to_pes_25_out_valid(PENetwork_9_io_to_pes_25_out_valid),
    .io_to_pes_25_out_bits(PENetwork_9_io_to_pes_25_out_bits),
    .io_to_pes_26_in_valid(PENetwork_9_io_to_pes_26_in_valid),
    .io_to_pes_26_in_bits(PENetwork_9_io_to_pes_26_in_bits),
    .io_to_pes_26_out_valid(PENetwork_9_io_to_pes_26_out_valid),
    .io_to_pes_26_out_bits(PENetwork_9_io_to_pes_26_out_bits),
    .io_to_pes_27_in_valid(PENetwork_9_io_to_pes_27_in_valid),
    .io_to_pes_27_in_bits(PENetwork_9_io_to_pes_27_in_bits),
    .io_to_pes_27_out_valid(PENetwork_9_io_to_pes_27_out_valid),
    .io_to_pes_27_out_bits(PENetwork_9_io_to_pes_27_out_bits),
    .io_to_pes_28_in_valid(PENetwork_9_io_to_pes_28_in_valid),
    .io_to_pes_28_in_bits(PENetwork_9_io_to_pes_28_in_bits),
    .io_to_pes_28_out_valid(PENetwork_9_io_to_pes_28_out_valid),
    .io_to_pes_28_out_bits(PENetwork_9_io_to_pes_28_out_bits),
    .io_to_pes_29_in_valid(PENetwork_9_io_to_pes_29_in_valid),
    .io_to_pes_29_in_bits(PENetwork_9_io_to_pes_29_in_bits),
    .io_to_mem_valid(PENetwork_9_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_9_io_to_mem_bits)
  );
  PENetwork PENetwork_10 ( // @[pe.scala 229:13]
    .io_to_pes_0_in_valid(PENetwork_10_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_10_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_10_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_10_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_10_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_10_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_10_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_10_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_10_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_10_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_10_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_10_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_10_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_10_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_10_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_10_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_10_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_10_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_10_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_10_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_10_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_10_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_10_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_10_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_10_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_10_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_10_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_10_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_10_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_10_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_10_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_10_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_10_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_10_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_10_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_10_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_10_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_10_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_10_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_10_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_10_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_10_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_10_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_10_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_10_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_10_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_10_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_10_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_10_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_10_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_10_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_10_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_10_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_10_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_10_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_10_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_10_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_10_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_10_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_10_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_10_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_10_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_10_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_10_io_to_pes_15_out_bits),
    .io_to_pes_16_in_valid(PENetwork_10_io_to_pes_16_in_valid),
    .io_to_pes_16_in_bits(PENetwork_10_io_to_pes_16_in_bits),
    .io_to_pes_16_out_valid(PENetwork_10_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_10_io_to_pes_16_out_bits),
    .io_to_pes_17_in_valid(PENetwork_10_io_to_pes_17_in_valid),
    .io_to_pes_17_in_bits(PENetwork_10_io_to_pes_17_in_bits),
    .io_to_pes_17_out_valid(PENetwork_10_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_10_io_to_pes_17_out_bits),
    .io_to_pes_18_in_valid(PENetwork_10_io_to_pes_18_in_valid),
    .io_to_pes_18_in_bits(PENetwork_10_io_to_pes_18_in_bits),
    .io_to_pes_18_out_valid(PENetwork_10_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_10_io_to_pes_18_out_bits),
    .io_to_pes_19_in_valid(PENetwork_10_io_to_pes_19_in_valid),
    .io_to_pes_19_in_bits(PENetwork_10_io_to_pes_19_in_bits),
    .io_to_pes_19_out_valid(PENetwork_10_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_10_io_to_pes_19_out_bits),
    .io_to_pes_20_in_valid(PENetwork_10_io_to_pes_20_in_valid),
    .io_to_pes_20_in_bits(PENetwork_10_io_to_pes_20_in_bits),
    .io_to_pes_20_out_valid(PENetwork_10_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_10_io_to_pes_20_out_bits),
    .io_to_pes_21_in_valid(PENetwork_10_io_to_pes_21_in_valid),
    .io_to_pes_21_in_bits(PENetwork_10_io_to_pes_21_in_bits),
    .io_to_pes_21_out_valid(PENetwork_10_io_to_pes_21_out_valid),
    .io_to_pes_21_out_bits(PENetwork_10_io_to_pes_21_out_bits),
    .io_to_pes_22_in_valid(PENetwork_10_io_to_pes_22_in_valid),
    .io_to_pes_22_in_bits(PENetwork_10_io_to_pes_22_in_bits),
    .io_to_pes_22_out_valid(PENetwork_10_io_to_pes_22_out_valid),
    .io_to_pes_22_out_bits(PENetwork_10_io_to_pes_22_out_bits),
    .io_to_pes_23_in_valid(PENetwork_10_io_to_pes_23_in_valid),
    .io_to_pes_23_in_bits(PENetwork_10_io_to_pes_23_in_bits),
    .io_to_pes_23_out_valid(PENetwork_10_io_to_pes_23_out_valid),
    .io_to_pes_23_out_bits(PENetwork_10_io_to_pes_23_out_bits),
    .io_to_pes_24_in_valid(PENetwork_10_io_to_pes_24_in_valid),
    .io_to_pes_24_in_bits(PENetwork_10_io_to_pes_24_in_bits),
    .io_to_pes_24_out_valid(PENetwork_10_io_to_pes_24_out_valid),
    .io_to_pes_24_out_bits(PENetwork_10_io_to_pes_24_out_bits),
    .io_to_pes_25_in_valid(PENetwork_10_io_to_pes_25_in_valid),
    .io_to_pes_25_in_bits(PENetwork_10_io_to_pes_25_in_bits),
    .io_to_pes_25_out_valid(PENetwork_10_io_to_pes_25_out_valid),
    .io_to_pes_25_out_bits(PENetwork_10_io_to_pes_25_out_bits),
    .io_to_pes_26_in_valid(PENetwork_10_io_to_pes_26_in_valid),
    .io_to_pes_26_in_bits(PENetwork_10_io_to_pes_26_in_bits),
    .io_to_pes_26_out_valid(PENetwork_10_io_to_pes_26_out_valid),
    .io_to_pes_26_out_bits(PENetwork_10_io_to_pes_26_out_bits),
    .io_to_pes_27_in_valid(PENetwork_10_io_to_pes_27_in_valid),
    .io_to_pes_27_in_bits(PENetwork_10_io_to_pes_27_in_bits),
    .io_to_pes_27_out_valid(PENetwork_10_io_to_pes_27_out_valid),
    .io_to_pes_27_out_bits(PENetwork_10_io_to_pes_27_out_bits),
    .io_to_pes_28_in_valid(PENetwork_10_io_to_pes_28_in_valid),
    .io_to_pes_28_in_bits(PENetwork_10_io_to_pes_28_in_bits),
    .io_to_pes_28_out_valid(PENetwork_10_io_to_pes_28_out_valid),
    .io_to_pes_28_out_bits(PENetwork_10_io_to_pes_28_out_bits),
    .io_to_pes_29_in_valid(PENetwork_10_io_to_pes_29_in_valid),
    .io_to_pes_29_in_bits(PENetwork_10_io_to_pes_29_in_bits),
    .io_to_mem_valid(PENetwork_10_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_10_io_to_mem_bits)
  );
  PENetwork PENetwork_11 ( // @[pe.scala 229:13]
    .io_to_pes_0_in_valid(PENetwork_11_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_11_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_11_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_11_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_11_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_11_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_11_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_11_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_11_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_11_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_11_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_11_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_11_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_11_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_11_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_11_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_11_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_11_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_11_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_11_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_11_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_11_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_11_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_11_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_11_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_11_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_11_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_11_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_11_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_11_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_11_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_11_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_11_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_11_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_11_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_11_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_11_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_11_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_11_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_11_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_11_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_11_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_11_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_11_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_11_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_11_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_11_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_11_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_11_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_11_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_11_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_11_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_11_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_11_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_11_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_11_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_11_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_11_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_11_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_11_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_11_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_11_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_11_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_11_io_to_pes_15_out_bits),
    .io_to_pes_16_in_valid(PENetwork_11_io_to_pes_16_in_valid),
    .io_to_pes_16_in_bits(PENetwork_11_io_to_pes_16_in_bits),
    .io_to_pes_16_out_valid(PENetwork_11_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_11_io_to_pes_16_out_bits),
    .io_to_pes_17_in_valid(PENetwork_11_io_to_pes_17_in_valid),
    .io_to_pes_17_in_bits(PENetwork_11_io_to_pes_17_in_bits),
    .io_to_pes_17_out_valid(PENetwork_11_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_11_io_to_pes_17_out_bits),
    .io_to_pes_18_in_valid(PENetwork_11_io_to_pes_18_in_valid),
    .io_to_pes_18_in_bits(PENetwork_11_io_to_pes_18_in_bits),
    .io_to_pes_18_out_valid(PENetwork_11_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_11_io_to_pes_18_out_bits),
    .io_to_pes_19_in_valid(PENetwork_11_io_to_pes_19_in_valid),
    .io_to_pes_19_in_bits(PENetwork_11_io_to_pes_19_in_bits),
    .io_to_pes_19_out_valid(PENetwork_11_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_11_io_to_pes_19_out_bits),
    .io_to_pes_20_in_valid(PENetwork_11_io_to_pes_20_in_valid),
    .io_to_pes_20_in_bits(PENetwork_11_io_to_pes_20_in_bits),
    .io_to_pes_20_out_valid(PENetwork_11_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_11_io_to_pes_20_out_bits),
    .io_to_pes_21_in_valid(PENetwork_11_io_to_pes_21_in_valid),
    .io_to_pes_21_in_bits(PENetwork_11_io_to_pes_21_in_bits),
    .io_to_pes_21_out_valid(PENetwork_11_io_to_pes_21_out_valid),
    .io_to_pes_21_out_bits(PENetwork_11_io_to_pes_21_out_bits),
    .io_to_pes_22_in_valid(PENetwork_11_io_to_pes_22_in_valid),
    .io_to_pes_22_in_bits(PENetwork_11_io_to_pes_22_in_bits),
    .io_to_pes_22_out_valid(PENetwork_11_io_to_pes_22_out_valid),
    .io_to_pes_22_out_bits(PENetwork_11_io_to_pes_22_out_bits),
    .io_to_pes_23_in_valid(PENetwork_11_io_to_pes_23_in_valid),
    .io_to_pes_23_in_bits(PENetwork_11_io_to_pes_23_in_bits),
    .io_to_pes_23_out_valid(PENetwork_11_io_to_pes_23_out_valid),
    .io_to_pes_23_out_bits(PENetwork_11_io_to_pes_23_out_bits),
    .io_to_pes_24_in_valid(PENetwork_11_io_to_pes_24_in_valid),
    .io_to_pes_24_in_bits(PENetwork_11_io_to_pes_24_in_bits),
    .io_to_pes_24_out_valid(PENetwork_11_io_to_pes_24_out_valid),
    .io_to_pes_24_out_bits(PENetwork_11_io_to_pes_24_out_bits),
    .io_to_pes_25_in_valid(PENetwork_11_io_to_pes_25_in_valid),
    .io_to_pes_25_in_bits(PENetwork_11_io_to_pes_25_in_bits),
    .io_to_pes_25_out_valid(PENetwork_11_io_to_pes_25_out_valid),
    .io_to_pes_25_out_bits(PENetwork_11_io_to_pes_25_out_bits),
    .io_to_pes_26_in_valid(PENetwork_11_io_to_pes_26_in_valid),
    .io_to_pes_26_in_bits(PENetwork_11_io_to_pes_26_in_bits),
    .io_to_pes_26_out_valid(PENetwork_11_io_to_pes_26_out_valid),
    .io_to_pes_26_out_bits(PENetwork_11_io_to_pes_26_out_bits),
    .io_to_pes_27_in_valid(PENetwork_11_io_to_pes_27_in_valid),
    .io_to_pes_27_in_bits(PENetwork_11_io_to_pes_27_in_bits),
    .io_to_pes_27_out_valid(PENetwork_11_io_to_pes_27_out_valid),
    .io_to_pes_27_out_bits(PENetwork_11_io_to_pes_27_out_bits),
    .io_to_pes_28_in_valid(PENetwork_11_io_to_pes_28_in_valid),
    .io_to_pes_28_in_bits(PENetwork_11_io_to_pes_28_in_bits),
    .io_to_pes_28_out_valid(PENetwork_11_io_to_pes_28_out_valid),
    .io_to_pes_28_out_bits(PENetwork_11_io_to_pes_28_out_bits),
    .io_to_pes_29_in_valid(PENetwork_11_io_to_pes_29_in_valid),
    .io_to_pes_29_in_bits(PENetwork_11_io_to_pes_29_in_bits),
    .io_to_mem_valid(PENetwork_11_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_11_io_to_mem_bits)
  );
  PENetwork PENetwork_12 ( // @[pe.scala 229:13]
    .io_to_pes_0_in_valid(PENetwork_12_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_12_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_12_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_12_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_12_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_12_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_12_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_12_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_12_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_12_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_12_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_12_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_12_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_12_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_12_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_12_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_12_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_12_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_12_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_12_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_12_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_12_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_12_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_12_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_12_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_12_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_12_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_12_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_12_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_12_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_12_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_12_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_12_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_12_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_12_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_12_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_12_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_12_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_12_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_12_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_12_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_12_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_12_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_12_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_12_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_12_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_12_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_12_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_12_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_12_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_12_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_12_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_12_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_12_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_12_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_12_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_12_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_12_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_12_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_12_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_12_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_12_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_12_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_12_io_to_pes_15_out_bits),
    .io_to_pes_16_in_valid(PENetwork_12_io_to_pes_16_in_valid),
    .io_to_pes_16_in_bits(PENetwork_12_io_to_pes_16_in_bits),
    .io_to_pes_16_out_valid(PENetwork_12_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_12_io_to_pes_16_out_bits),
    .io_to_pes_17_in_valid(PENetwork_12_io_to_pes_17_in_valid),
    .io_to_pes_17_in_bits(PENetwork_12_io_to_pes_17_in_bits),
    .io_to_pes_17_out_valid(PENetwork_12_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_12_io_to_pes_17_out_bits),
    .io_to_pes_18_in_valid(PENetwork_12_io_to_pes_18_in_valid),
    .io_to_pes_18_in_bits(PENetwork_12_io_to_pes_18_in_bits),
    .io_to_pes_18_out_valid(PENetwork_12_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_12_io_to_pes_18_out_bits),
    .io_to_pes_19_in_valid(PENetwork_12_io_to_pes_19_in_valid),
    .io_to_pes_19_in_bits(PENetwork_12_io_to_pes_19_in_bits),
    .io_to_pes_19_out_valid(PENetwork_12_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_12_io_to_pes_19_out_bits),
    .io_to_pes_20_in_valid(PENetwork_12_io_to_pes_20_in_valid),
    .io_to_pes_20_in_bits(PENetwork_12_io_to_pes_20_in_bits),
    .io_to_pes_20_out_valid(PENetwork_12_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_12_io_to_pes_20_out_bits),
    .io_to_pes_21_in_valid(PENetwork_12_io_to_pes_21_in_valid),
    .io_to_pes_21_in_bits(PENetwork_12_io_to_pes_21_in_bits),
    .io_to_pes_21_out_valid(PENetwork_12_io_to_pes_21_out_valid),
    .io_to_pes_21_out_bits(PENetwork_12_io_to_pes_21_out_bits),
    .io_to_pes_22_in_valid(PENetwork_12_io_to_pes_22_in_valid),
    .io_to_pes_22_in_bits(PENetwork_12_io_to_pes_22_in_bits),
    .io_to_pes_22_out_valid(PENetwork_12_io_to_pes_22_out_valid),
    .io_to_pes_22_out_bits(PENetwork_12_io_to_pes_22_out_bits),
    .io_to_pes_23_in_valid(PENetwork_12_io_to_pes_23_in_valid),
    .io_to_pes_23_in_bits(PENetwork_12_io_to_pes_23_in_bits),
    .io_to_pes_23_out_valid(PENetwork_12_io_to_pes_23_out_valid),
    .io_to_pes_23_out_bits(PENetwork_12_io_to_pes_23_out_bits),
    .io_to_pes_24_in_valid(PENetwork_12_io_to_pes_24_in_valid),
    .io_to_pes_24_in_bits(PENetwork_12_io_to_pes_24_in_bits),
    .io_to_pes_24_out_valid(PENetwork_12_io_to_pes_24_out_valid),
    .io_to_pes_24_out_bits(PENetwork_12_io_to_pes_24_out_bits),
    .io_to_pes_25_in_valid(PENetwork_12_io_to_pes_25_in_valid),
    .io_to_pes_25_in_bits(PENetwork_12_io_to_pes_25_in_bits),
    .io_to_pes_25_out_valid(PENetwork_12_io_to_pes_25_out_valid),
    .io_to_pes_25_out_bits(PENetwork_12_io_to_pes_25_out_bits),
    .io_to_pes_26_in_valid(PENetwork_12_io_to_pes_26_in_valid),
    .io_to_pes_26_in_bits(PENetwork_12_io_to_pes_26_in_bits),
    .io_to_pes_26_out_valid(PENetwork_12_io_to_pes_26_out_valid),
    .io_to_pes_26_out_bits(PENetwork_12_io_to_pes_26_out_bits),
    .io_to_pes_27_in_valid(PENetwork_12_io_to_pes_27_in_valid),
    .io_to_pes_27_in_bits(PENetwork_12_io_to_pes_27_in_bits),
    .io_to_pes_27_out_valid(PENetwork_12_io_to_pes_27_out_valid),
    .io_to_pes_27_out_bits(PENetwork_12_io_to_pes_27_out_bits),
    .io_to_pes_28_in_valid(PENetwork_12_io_to_pes_28_in_valid),
    .io_to_pes_28_in_bits(PENetwork_12_io_to_pes_28_in_bits),
    .io_to_pes_28_out_valid(PENetwork_12_io_to_pes_28_out_valid),
    .io_to_pes_28_out_bits(PENetwork_12_io_to_pes_28_out_bits),
    .io_to_pes_29_in_valid(PENetwork_12_io_to_pes_29_in_valid),
    .io_to_pes_29_in_bits(PENetwork_12_io_to_pes_29_in_bits),
    .io_to_mem_valid(PENetwork_12_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_12_io_to_mem_bits)
  );
  PENetwork PENetwork_13 ( // @[pe.scala 229:13]
    .io_to_pes_0_in_valid(PENetwork_13_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_13_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_13_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_13_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_13_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_13_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_13_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_13_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_13_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_13_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_13_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_13_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_13_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_13_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_13_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_13_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_13_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_13_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_13_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_13_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_13_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_13_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_13_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_13_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_13_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_13_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_13_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_13_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_13_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_13_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_13_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_13_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_13_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_13_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_13_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_13_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_13_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_13_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_13_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_13_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_13_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_13_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_13_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_13_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_13_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_13_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_13_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_13_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_13_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_13_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_13_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_13_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_13_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_13_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_13_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_13_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_13_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_13_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_13_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_13_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_13_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_13_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_13_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_13_io_to_pes_15_out_bits),
    .io_to_pes_16_in_valid(PENetwork_13_io_to_pes_16_in_valid),
    .io_to_pes_16_in_bits(PENetwork_13_io_to_pes_16_in_bits),
    .io_to_pes_16_out_valid(PENetwork_13_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_13_io_to_pes_16_out_bits),
    .io_to_pes_17_in_valid(PENetwork_13_io_to_pes_17_in_valid),
    .io_to_pes_17_in_bits(PENetwork_13_io_to_pes_17_in_bits),
    .io_to_pes_17_out_valid(PENetwork_13_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_13_io_to_pes_17_out_bits),
    .io_to_pes_18_in_valid(PENetwork_13_io_to_pes_18_in_valid),
    .io_to_pes_18_in_bits(PENetwork_13_io_to_pes_18_in_bits),
    .io_to_pes_18_out_valid(PENetwork_13_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_13_io_to_pes_18_out_bits),
    .io_to_pes_19_in_valid(PENetwork_13_io_to_pes_19_in_valid),
    .io_to_pes_19_in_bits(PENetwork_13_io_to_pes_19_in_bits),
    .io_to_pes_19_out_valid(PENetwork_13_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_13_io_to_pes_19_out_bits),
    .io_to_pes_20_in_valid(PENetwork_13_io_to_pes_20_in_valid),
    .io_to_pes_20_in_bits(PENetwork_13_io_to_pes_20_in_bits),
    .io_to_pes_20_out_valid(PENetwork_13_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_13_io_to_pes_20_out_bits),
    .io_to_pes_21_in_valid(PENetwork_13_io_to_pes_21_in_valid),
    .io_to_pes_21_in_bits(PENetwork_13_io_to_pes_21_in_bits),
    .io_to_pes_21_out_valid(PENetwork_13_io_to_pes_21_out_valid),
    .io_to_pes_21_out_bits(PENetwork_13_io_to_pes_21_out_bits),
    .io_to_pes_22_in_valid(PENetwork_13_io_to_pes_22_in_valid),
    .io_to_pes_22_in_bits(PENetwork_13_io_to_pes_22_in_bits),
    .io_to_pes_22_out_valid(PENetwork_13_io_to_pes_22_out_valid),
    .io_to_pes_22_out_bits(PENetwork_13_io_to_pes_22_out_bits),
    .io_to_pes_23_in_valid(PENetwork_13_io_to_pes_23_in_valid),
    .io_to_pes_23_in_bits(PENetwork_13_io_to_pes_23_in_bits),
    .io_to_pes_23_out_valid(PENetwork_13_io_to_pes_23_out_valid),
    .io_to_pes_23_out_bits(PENetwork_13_io_to_pes_23_out_bits),
    .io_to_pes_24_in_valid(PENetwork_13_io_to_pes_24_in_valid),
    .io_to_pes_24_in_bits(PENetwork_13_io_to_pes_24_in_bits),
    .io_to_pes_24_out_valid(PENetwork_13_io_to_pes_24_out_valid),
    .io_to_pes_24_out_bits(PENetwork_13_io_to_pes_24_out_bits),
    .io_to_pes_25_in_valid(PENetwork_13_io_to_pes_25_in_valid),
    .io_to_pes_25_in_bits(PENetwork_13_io_to_pes_25_in_bits),
    .io_to_pes_25_out_valid(PENetwork_13_io_to_pes_25_out_valid),
    .io_to_pes_25_out_bits(PENetwork_13_io_to_pes_25_out_bits),
    .io_to_pes_26_in_valid(PENetwork_13_io_to_pes_26_in_valid),
    .io_to_pes_26_in_bits(PENetwork_13_io_to_pes_26_in_bits),
    .io_to_pes_26_out_valid(PENetwork_13_io_to_pes_26_out_valid),
    .io_to_pes_26_out_bits(PENetwork_13_io_to_pes_26_out_bits),
    .io_to_pes_27_in_valid(PENetwork_13_io_to_pes_27_in_valid),
    .io_to_pes_27_in_bits(PENetwork_13_io_to_pes_27_in_bits),
    .io_to_pes_27_out_valid(PENetwork_13_io_to_pes_27_out_valid),
    .io_to_pes_27_out_bits(PENetwork_13_io_to_pes_27_out_bits),
    .io_to_pes_28_in_valid(PENetwork_13_io_to_pes_28_in_valid),
    .io_to_pes_28_in_bits(PENetwork_13_io_to_pes_28_in_bits),
    .io_to_pes_28_out_valid(PENetwork_13_io_to_pes_28_out_valid),
    .io_to_pes_28_out_bits(PENetwork_13_io_to_pes_28_out_bits),
    .io_to_pes_29_in_valid(PENetwork_13_io_to_pes_29_in_valid),
    .io_to_pes_29_in_bits(PENetwork_13_io_to_pes_29_in_bits),
    .io_to_mem_valid(PENetwork_13_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_13_io_to_mem_bits)
  );
  PENetwork PENetwork_14 ( // @[pe.scala 229:13]
    .io_to_pes_0_in_valid(PENetwork_14_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_14_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_14_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_14_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_14_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_14_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_14_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_14_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_14_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_14_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_14_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_14_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_14_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_14_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_14_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_14_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_14_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_14_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_14_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_14_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_14_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_14_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_14_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_14_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_14_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_14_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_14_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_14_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_14_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_14_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_14_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_14_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_14_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_14_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_14_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_14_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_14_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_14_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_14_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_14_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_14_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_14_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_14_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_14_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_14_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_14_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_14_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_14_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_14_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_14_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_14_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_14_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_14_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_14_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_14_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_14_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_14_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_14_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_14_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_14_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_14_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_14_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_14_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_14_io_to_pes_15_out_bits),
    .io_to_pes_16_in_valid(PENetwork_14_io_to_pes_16_in_valid),
    .io_to_pes_16_in_bits(PENetwork_14_io_to_pes_16_in_bits),
    .io_to_pes_16_out_valid(PENetwork_14_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_14_io_to_pes_16_out_bits),
    .io_to_pes_17_in_valid(PENetwork_14_io_to_pes_17_in_valid),
    .io_to_pes_17_in_bits(PENetwork_14_io_to_pes_17_in_bits),
    .io_to_pes_17_out_valid(PENetwork_14_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_14_io_to_pes_17_out_bits),
    .io_to_pes_18_in_valid(PENetwork_14_io_to_pes_18_in_valid),
    .io_to_pes_18_in_bits(PENetwork_14_io_to_pes_18_in_bits),
    .io_to_pes_18_out_valid(PENetwork_14_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_14_io_to_pes_18_out_bits),
    .io_to_pes_19_in_valid(PENetwork_14_io_to_pes_19_in_valid),
    .io_to_pes_19_in_bits(PENetwork_14_io_to_pes_19_in_bits),
    .io_to_pes_19_out_valid(PENetwork_14_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_14_io_to_pes_19_out_bits),
    .io_to_pes_20_in_valid(PENetwork_14_io_to_pes_20_in_valid),
    .io_to_pes_20_in_bits(PENetwork_14_io_to_pes_20_in_bits),
    .io_to_pes_20_out_valid(PENetwork_14_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_14_io_to_pes_20_out_bits),
    .io_to_pes_21_in_valid(PENetwork_14_io_to_pes_21_in_valid),
    .io_to_pes_21_in_bits(PENetwork_14_io_to_pes_21_in_bits),
    .io_to_pes_21_out_valid(PENetwork_14_io_to_pes_21_out_valid),
    .io_to_pes_21_out_bits(PENetwork_14_io_to_pes_21_out_bits),
    .io_to_pes_22_in_valid(PENetwork_14_io_to_pes_22_in_valid),
    .io_to_pes_22_in_bits(PENetwork_14_io_to_pes_22_in_bits),
    .io_to_pes_22_out_valid(PENetwork_14_io_to_pes_22_out_valid),
    .io_to_pes_22_out_bits(PENetwork_14_io_to_pes_22_out_bits),
    .io_to_pes_23_in_valid(PENetwork_14_io_to_pes_23_in_valid),
    .io_to_pes_23_in_bits(PENetwork_14_io_to_pes_23_in_bits),
    .io_to_pes_23_out_valid(PENetwork_14_io_to_pes_23_out_valid),
    .io_to_pes_23_out_bits(PENetwork_14_io_to_pes_23_out_bits),
    .io_to_pes_24_in_valid(PENetwork_14_io_to_pes_24_in_valid),
    .io_to_pes_24_in_bits(PENetwork_14_io_to_pes_24_in_bits),
    .io_to_pes_24_out_valid(PENetwork_14_io_to_pes_24_out_valid),
    .io_to_pes_24_out_bits(PENetwork_14_io_to_pes_24_out_bits),
    .io_to_pes_25_in_valid(PENetwork_14_io_to_pes_25_in_valid),
    .io_to_pes_25_in_bits(PENetwork_14_io_to_pes_25_in_bits),
    .io_to_pes_25_out_valid(PENetwork_14_io_to_pes_25_out_valid),
    .io_to_pes_25_out_bits(PENetwork_14_io_to_pes_25_out_bits),
    .io_to_pes_26_in_valid(PENetwork_14_io_to_pes_26_in_valid),
    .io_to_pes_26_in_bits(PENetwork_14_io_to_pes_26_in_bits),
    .io_to_pes_26_out_valid(PENetwork_14_io_to_pes_26_out_valid),
    .io_to_pes_26_out_bits(PENetwork_14_io_to_pes_26_out_bits),
    .io_to_pes_27_in_valid(PENetwork_14_io_to_pes_27_in_valid),
    .io_to_pes_27_in_bits(PENetwork_14_io_to_pes_27_in_bits),
    .io_to_pes_27_out_valid(PENetwork_14_io_to_pes_27_out_valid),
    .io_to_pes_27_out_bits(PENetwork_14_io_to_pes_27_out_bits),
    .io_to_pes_28_in_valid(PENetwork_14_io_to_pes_28_in_valid),
    .io_to_pes_28_in_bits(PENetwork_14_io_to_pes_28_in_bits),
    .io_to_pes_28_out_valid(PENetwork_14_io_to_pes_28_out_valid),
    .io_to_pes_28_out_bits(PENetwork_14_io_to_pes_28_out_bits),
    .io_to_pes_29_in_valid(PENetwork_14_io_to_pes_29_in_valid),
    .io_to_pes_29_in_bits(PENetwork_14_io_to_pes_29_in_bits),
    .io_to_mem_valid(PENetwork_14_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_14_io_to_mem_bits)
  );
  PENetwork PENetwork_15 ( // @[pe.scala 229:13]
    .io_to_pes_0_in_valid(PENetwork_15_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_15_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_15_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_15_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_15_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_15_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_15_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_15_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_15_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_15_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_15_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_15_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_15_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_15_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_15_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_15_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_15_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_15_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_15_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_15_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_15_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_15_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_15_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_15_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_15_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_15_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_15_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_15_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_15_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_15_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_15_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_15_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_15_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_15_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_15_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_15_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_15_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_15_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_15_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_15_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_15_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_15_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_15_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_15_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_15_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_15_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_15_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_15_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_15_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_15_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_15_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_15_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_15_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_15_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_15_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_15_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_15_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_15_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_15_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_15_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_15_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_15_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_15_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_15_io_to_pes_15_out_bits),
    .io_to_pes_16_in_valid(PENetwork_15_io_to_pes_16_in_valid),
    .io_to_pes_16_in_bits(PENetwork_15_io_to_pes_16_in_bits),
    .io_to_pes_16_out_valid(PENetwork_15_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_15_io_to_pes_16_out_bits),
    .io_to_pes_17_in_valid(PENetwork_15_io_to_pes_17_in_valid),
    .io_to_pes_17_in_bits(PENetwork_15_io_to_pes_17_in_bits),
    .io_to_pes_17_out_valid(PENetwork_15_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_15_io_to_pes_17_out_bits),
    .io_to_pes_18_in_valid(PENetwork_15_io_to_pes_18_in_valid),
    .io_to_pes_18_in_bits(PENetwork_15_io_to_pes_18_in_bits),
    .io_to_pes_18_out_valid(PENetwork_15_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_15_io_to_pes_18_out_bits),
    .io_to_pes_19_in_valid(PENetwork_15_io_to_pes_19_in_valid),
    .io_to_pes_19_in_bits(PENetwork_15_io_to_pes_19_in_bits),
    .io_to_pes_19_out_valid(PENetwork_15_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_15_io_to_pes_19_out_bits),
    .io_to_pes_20_in_valid(PENetwork_15_io_to_pes_20_in_valid),
    .io_to_pes_20_in_bits(PENetwork_15_io_to_pes_20_in_bits),
    .io_to_pes_20_out_valid(PENetwork_15_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_15_io_to_pes_20_out_bits),
    .io_to_pes_21_in_valid(PENetwork_15_io_to_pes_21_in_valid),
    .io_to_pes_21_in_bits(PENetwork_15_io_to_pes_21_in_bits),
    .io_to_pes_21_out_valid(PENetwork_15_io_to_pes_21_out_valid),
    .io_to_pes_21_out_bits(PENetwork_15_io_to_pes_21_out_bits),
    .io_to_pes_22_in_valid(PENetwork_15_io_to_pes_22_in_valid),
    .io_to_pes_22_in_bits(PENetwork_15_io_to_pes_22_in_bits),
    .io_to_pes_22_out_valid(PENetwork_15_io_to_pes_22_out_valid),
    .io_to_pes_22_out_bits(PENetwork_15_io_to_pes_22_out_bits),
    .io_to_pes_23_in_valid(PENetwork_15_io_to_pes_23_in_valid),
    .io_to_pes_23_in_bits(PENetwork_15_io_to_pes_23_in_bits),
    .io_to_pes_23_out_valid(PENetwork_15_io_to_pes_23_out_valid),
    .io_to_pes_23_out_bits(PENetwork_15_io_to_pes_23_out_bits),
    .io_to_pes_24_in_valid(PENetwork_15_io_to_pes_24_in_valid),
    .io_to_pes_24_in_bits(PENetwork_15_io_to_pes_24_in_bits),
    .io_to_pes_24_out_valid(PENetwork_15_io_to_pes_24_out_valid),
    .io_to_pes_24_out_bits(PENetwork_15_io_to_pes_24_out_bits),
    .io_to_pes_25_in_valid(PENetwork_15_io_to_pes_25_in_valid),
    .io_to_pes_25_in_bits(PENetwork_15_io_to_pes_25_in_bits),
    .io_to_pes_25_out_valid(PENetwork_15_io_to_pes_25_out_valid),
    .io_to_pes_25_out_bits(PENetwork_15_io_to_pes_25_out_bits),
    .io_to_pes_26_in_valid(PENetwork_15_io_to_pes_26_in_valid),
    .io_to_pes_26_in_bits(PENetwork_15_io_to_pes_26_in_bits),
    .io_to_pes_26_out_valid(PENetwork_15_io_to_pes_26_out_valid),
    .io_to_pes_26_out_bits(PENetwork_15_io_to_pes_26_out_bits),
    .io_to_pes_27_in_valid(PENetwork_15_io_to_pes_27_in_valid),
    .io_to_pes_27_in_bits(PENetwork_15_io_to_pes_27_in_bits),
    .io_to_pes_27_out_valid(PENetwork_15_io_to_pes_27_out_valid),
    .io_to_pes_27_out_bits(PENetwork_15_io_to_pes_27_out_bits),
    .io_to_pes_28_in_valid(PENetwork_15_io_to_pes_28_in_valid),
    .io_to_pes_28_in_bits(PENetwork_15_io_to_pes_28_in_bits),
    .io_to_pes_28_out_valid(PENetwork_15_io_to_pes_28_out_valid),
    .io_to_pes_28_out_bits(PENetwork_15_io_to_pes_28_out_bits),
    .io_to_pes_29_in_valid(PENetwork_15_io_to_pes_29_in_valid),
    .io_to_pes_29_in_bits(PENetwork_15_io_to_pes_29_in_bits),
    .io_to_mem_valid(PENetwork_15_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_15_io_to_mem_bits)
  );
  PENetwork PENetwork_16 ( // @[pe.scala 229:13]
    .io_to_pes_0_in_valid(PENetwork_16_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_16_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_16_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_16_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_16_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_16_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_16_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_16_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_16_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_16_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_16_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_16_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_16_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_16_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_16_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_16_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_16_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_16_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_16_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_16_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_16_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_16_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_16_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_16_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_16_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_16_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_16_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_16_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_16_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_16_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_16_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_16_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_16_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_16_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_16_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_16_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_16_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_16_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_16_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_16_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_16_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_16_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_16_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_16_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_16_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_16_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_16_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_16_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_16_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_16_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_16_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_16_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_16_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_16_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_16_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_16_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_16_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_16_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_16_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_16_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_16_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_16_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_16_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_16_io_to_pes_15_out_bits),
    .io_to_pes_16_in_valid(PENetwork_16_io_to_pes_16_in_valid),
    .io_to_pes_16_in_bits(PENetwork_16_io_to_pes_16_in_bits),
    .io_to_pes_16_out_valid(PENetwork_16_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_16_io_to_pes_16_out_bits),
    .io_to_pes_17_in_valid(PENetwork_16_io_to_pes_17_in_valid),
    .io_to_pes_17_in_bits(PENetwork_16_io_to_pes_17_in_bits),
    .io_to_pes_17_out_valid(PENetwork_16_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_16_io_to_pes_17_out_bits),
    .io_to_pes_18_in_valid(PENetwork_16_io_to_pes_18_in_valid),
    .io_to_pes_18_in_bits(PENetwork_16_io_to_pes_18_in_bits),
    .io_to_pes_18_out_valid(PENetwork_16_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_16_io_to_pes_18_out_bits),
    .io_to_pes_19_in_valid(PENetwork_16_io_to_pes_19_in_valid),
    .io_to_pes_19_in_bits(PENetwork_16_io_to_pes_19_in_bits),
    .io_to_pes_19_out_valid(PENetwork_16_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_16_io_to_pes_19_out_bits),
    .io_to_pes_20_in_valid(PENetwork_16_io_to_pes_20_in_valid),
    .io_to_pes_20_in_bits(PENetwork_16_io_to_pes_20_in_bits),
    .io_to_pes_20_out_valid(PENetwork_16_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_16_io_to_pes_20_out_bits),
    .io_to_pes_21_in_valid(PENetwork_16_io_to_pes_21_in_valid),
    .io_to_pes_21_in_bits(PENetwork_16_io_to_pes_21_in_bits),
    .io_to_pes_21_out_valid(PENetwork_16_io_to_pes_21_out_valid),
    .io_to_pes_21_out_bits(PENetwork_16_io_to_pes_21_out_bits),
    .io_to_pes_22_in_valid(PENetwork_16_io_to_pes_22_in_valid),
    .io_to_pes_22_in_bits(PENetwork_16_io_to_pes_22_in_bits),
    .io_to_pes_22_out_valid(PENetwork_16_io_to_pes_22_out_valid),
    .io_to_pes_22_out_bits(PENetwork_16_io_to_pes_22_out_bits),
    .io_to_pes_23_in_valid(PENetwork_16_io_to_pes_23_in_valid),
    .io_to_pes_23_in_bits(PENetwork_16_io_to_pes_23_in_bits),
    .io_to_pes_23_out_valid(PENetwork_16_io_to_pes_23_out_valid),
    .io_to_pes_23_out_bits(PENetwork_16_io_to_pes_23_out_bits),
    .io_to_pes_24_in_valid(PENetwork_16_io_to_pes_24_in_valid),
    .io_to_pes_24_in_bits(PENetwork_16_io_to_pes_24_in_bits),
    .io_to_pes_24_out_valid(PENetwork_16_io_to_pes_24_out_valid),
    .io_to_pes_24_out_bits(PENetwork_16_io_to_pes_24_out_bits),
    .io_to_pes_25_in_valid(PENetwork_16_io_to_pes_25_in_valid),
    .io_to_pes_25_in_bits(PENetwork_16_io_to_pes_25_in_bits),
    .io_to_pes_25_out_valid(PENetwork_16_io_to_pes_25_out_valid),
    .io_to_pes_25_out_bits(PENetwork_16_io_to_pes_25_out_bits),
    .io_to_pes_26_in_valid(PENetwork_16_io_to_pes_26_in_valid),
    .io_to_pes_26_in_bits(PENetwork_16_io_to_pes_26_in_bits),
    .io_to_pes_26_out_valid(PENetwork_16_io_to_pes_26_out_valid),
    .io_to_pes_26_out_bits(PENetwork_16_io_to_pes_26_out_bits),
    .io_to_pes_27_in_valid(PENetwork_16_io_to_pes_27_in_valid),
    .io_to_pes_27_in_bits(PENetwork_16_io_to_pes_27_in_bits),
    .io_to_pes_27_out_valid(PENetwork_16_io_to_pes_27_out_valid),
    .io_to_pes_27_out_bits(PENetwork_16_io_to_pes_27_out_bits),
    .io_to_pes_28_in_valid(PENetwork_16_io_to_pes_28_in_valid),
    .io_to_pes_28_in_bits(PENetwork_16_io_to_pes_28_in_bits),
    .io_to_pes_28_out_valid(PENetwork_16_io_to_pes_28_out_valid),
    .io_to_pes_28_out_bits(PENetwork_16_io_to_pes_28_out_bits),
    .io_to_pes_29_in_valid(PENetwork_16_io_to_pes_29_in_valid),
    .io_to_pes_29_in_bits(PENetwork_16_io_to_pes_29_in_bits),
    .io_to_mem_valid(PENetwork_16_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_16_io_to_mem_bits)
  );
  PENetwork PENetwork_17 ( // @[pe.scala 229:13]
    .io_to_pes_0_in_valid(PENetwork_17_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_17_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_17_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_17_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_17_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_17_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_17_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_17_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_17_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_17_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_17_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_17_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_17_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_17_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_17_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_17_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_17_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_17_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_17_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_17_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_17_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_17_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_17_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_17_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_17_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_17_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_17_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_17_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_17_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_17_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_17_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_17_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_17_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_17_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_17_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_17_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_17_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_17_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_17_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_17_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_17_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_17_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_17_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_17_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_17_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_17_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_17_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_17_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_17_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_17_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_17_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_17_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_17_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_17_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_17_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_17_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_17_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_17_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_17_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_17_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_17_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_17_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_17_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_17_io_to_pes_15_out_bits),
    .io_to_pes_16_in_valid(PENetwork_17_io_to_pes_16_in_valid),
    .io_to_pes_16_in_bits(PENetwork_17_io_to_pes_16_in_bits),
    .io_to_pes_16_out_valid(PENetwork_17_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_17_io_to_pes_16_out_bits),
    .io_to_pes_17_in_valid(PENetwork_17_io_to_pes_17_in_valid),
    .io_to_pes_17_in_bits(PENetwork_17_io_to_pes_17_in_bits),
    .io_to_pes_17_out_valid(PENetwork_17_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_17_io_to_pes_17_out_bits),
    .io_to_pes_18_in_valid(PENetwork_17_io_to_pes_18_in_valid),
    .io_to_pes_18_in_bits(PENetwork_17_io_to_pes_18_in_bits),
    .io_to_pes_18_out_valid(PENetwork_17_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_17_io_to_pes_18_out_bits),
    .io_to_pes_19_in_valid(PENetwork_17_io_to_pes_19_in_valid),
    .io_to_pes_19_in_bits(PENetwork_17_io_to_pes_19_in_bits),
    .io_to_pes_19_out_valid(PENetwork_17_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_17_io_to_pes_19_out_bits),
    .io_to_pes_20_in_valid(PENetwork_17_io_to_pes_20_in_valid),
    .io_to_pes_20_in_bits(PENetwork_17_io_to_pes_20_in_bits),
    .io_to_pes_20_out_valid(PENetwork_17_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_17_io_to_pes_20_out_bits),
    .io_to_pes_21_in_valid(PENetwork_17_io_to_pes_21_in_valid),
    .io_to_pes_21_in_bits(PENetwork_17_io_to_pes_21_in_bits),
    .io_to_pes_21_out_valid(PENetwork_17_io_to_pes_21_out_valid),
    .io_to_pes_21_out_bits(PENetwork_17_io_to_pes_21_out_bits),
    .io_to_pes_22_in_valid(PENetwork_17_io_to_pes_22_in_valid),
    .io_to_pes_22_in_bits(PENetwork_17_io_to_pes_22_in_bits),
    .io_to_pes_22_out_valid(PENetwork_17_io_to_pes_22_out_valid),
    .io_to_pes_22_out_bits(PENetwork_17_io_to_pes_22_out_bits),
    .io_to_pes_23_in_valid(PENetwork_17_io_to_pes_23_in_valid),
    .io_to_pes_23_in_bits(PENetwork_17_io_to_pes_23_in_bits),
    .io_to_pes_23_out_valid(PENetwork_17_io_to_pes_23_out_valid),
    .io_to_pes_23_out_bits(PENetwork_17_io_to_pes_23_out_bits),
    .io_to_pes_24_in_valid(PENetwork_17_io_to_pes_24_in_valid),
    .io_to_pes_24_in_bits(PENetwork_17_io_to_pes_24_in_bits),
    .io_to_pes_24_out_valid(PENetwork_17_io_to_pes_24_out_valid),
    .io_to_pes_24_out_bits(PENetwork_17_io_to_pes_24_out_bits),
    .io_to_pes_25_in_valid(PENetwork_17_io_to_pes_25_in_valid),
    .io_to_pes_25_in_bits(PENetwork_17_io_to_pes_25_in_bits),
    .io_to_pes_25_out_valid(PENetwork_17_io_to_pes_25_out_valid),
    .io_to_pes_25_out_bits(PENetwork_17_io_to_pes_25_out_bits),
    .io_to_pes_26_in_valid(PENetwork_17_io_to_pes_26_in_valid),
    .io_to_pes_26_in_bits(PENetwork_17_io_to_pes_26_in_bits),
    .io_to_pes_26_out_valid(PENetwork_17_io_to_pes_26_out_valid),
    .io_to_pes_26_out_bits(PENetwork_17_io_to_pes_26_out_bits),
    .io_to_pes_27_in_valid(PENetwork_17_io_to_pes_27_in_valid),
    .io_to_pes_27_in_bits(PENetwork_17_io_to_pes_27_in_bits),
    .io_to_pes_27_out_valid(PENetwork_17_io_to_pes_27_out_valid),
    .io_to_pes_27_out_bits(PENetwork_17_io_to_pes_27_out_bits),
    .io_to_pes_28_in_valid(PENetwork_17_io_to_pes_28_in_valid),
    .io_to_pes_28_in_bits(PENetwork_17_io_to_pes_28_in_bits),
    .io_to_pes_28_out_valid(PENetwork_17_io_to_pes_28_out_valid),
    .io_to_pes_28_out_bits(PENetwork_17_io_to_pes_28_out_bits),
    .io_to_pes_29_in_valid(PENetwork_17_io_to_pes_29_in_valid),
    .io_to_pes_29_in_bits(PENetwork_17_io_to_pes_29_in_bits),
    .io_to_mem_valid(PENetwork_17_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_17_io_to_mem_bits)
  );
  PENetwork PENetwork_18 ( // @[pe.scala 229:13]
    .io_to_pes_0_in_valid(PENetwork_18_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_18_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_18_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_18_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_18_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_18_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_18_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_18_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_18_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_18_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_18_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_18_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_18_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_18_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_18_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_18_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_18_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_18_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_18_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_18_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_18_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_18_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_18_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_18_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_18_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_18_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_18_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_18_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_18_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_18_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_18_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_18_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_18_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_18_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_18_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_18_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_18_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_18_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_18_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_18_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_18_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_18_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_18_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_18_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_18_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_18_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_18_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_18_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_18_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_18_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_18_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_18_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_18_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_18_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_18_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_18_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_18_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_18_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_18_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_18_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_18_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_18_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_18_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_18_io_to_pes_15_out_bits),
    .io_to_pes_16_in_valid(PENetwork_18_io_to_pes_16_in_valid),
    .io_to_pes_16_in_bits(PENetwork_18_io_to_pes_16_in_bits),
    .io_to_pes_16_out_valid(PENetwork_18_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_18_io_to_pes_16_out_bits),
    .io_to_pes_17_in_valid(PENetwork_18_io_to_pes_17_in_valid),
    .io_to_pes_17_in_bits(PENetwork_18_io_to_pes_17_in_bits),
    .io_to_pes_17_out_valid(PENetwork_18_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_18_io_to_pes_17_out_bits),
    .io_to_pes_18_in_valid(PENetwork_18_io_to_pes_18_in_valid),
    .io_to_pes_18_in_bits(PENetwork_18_io_to_pes_18_in_bits),
    .io_to_pes_18_out_valid(PENetwork_18_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_18_io_to_pes_18_out_bits),
    .io_to_pes_19_in_valid(PENetwork_18_io_to_pes_19_in_valid),
    .io_to_pes_19_in_bits(PENetwork_18_io_to_pes_19_in_bits),
    .io_to_pes_19_out_valid(PENetwork_18_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_18_io_to_pes_19_out_bits),
    .io_to_pes_20_in_valid(PENetwork_18_io_to_pes_20_in_valid),
    .io_to_pes_20_in_bits(PENetwork_18_io_to_pes_20_in_bits),
    .io_to_pes_20_out_valid(PENetwork_18_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_18_io_to_pes_20_out_bits),
    .io_to_pes_21_in_valid(PENetwork_18_io_to_pes_21_in_valid),
    .io_to_pes_21_in_bits(PENetwork_18_io_to_pes_21_in_bits),
    .io_to_pes_21_out_valid(PENetwork_18_io_to_pes_21_out_valid),
    .io_to_pes_21_out_bits(PENetwork_18_io_to_pes_21_out_bits),
    .io_to_pes_22_in_valid(PENetwork_18_io_to_pes_22_in_valid),
    .io_to_pes_22_in_bits(PENetwork_18_io_to_pes_22_in_bits),
    .io_to_pes_22_out_valid(PENetwork_18_io_to_pes_22_out_valid),
    .io_to_pes_22_out_bits(PENetwork_18_io_to_pes_22_out_bits),
    .io_to_pes_23_in_valid(PENetwork_18_io_to_pes_23_in_valid),
    .io_to_pes_23_in_bits(PENetwork_18_io_to_pes_23_in_bits),
    .io_to_pes_23_out_valid(PENetwork_18_io_to_pes_23_out_valid),
    .io_to_pes_23_out_bits(PENetwork_18_io_to_pes_23_out_bits),
    .io_to_pes_24_in_valid(PENetwork_18_io_to_pes_24_in_valid),
    .io_to_pes_24_in_bits(PENetwork_18_io_to_pes_24_in_bits),
    .io_to_pes_24_out_valid(PENetwork_18_io_to_pes_24_out_valid),
    .io_to_pes_24_out_bits(PENetwork_18_io_to_pes_24_out_bits),
    .io_to_pes_25_in_valid(PENetwork_18_io_to_pes_25_in_valid),
    .io_to_pes_25_in_bits(PENetwork_18_io_to_pes_25_in_bits),
    .io_to_pes_25_out_valid(PENetwork_18_io_to_pes_25_out_valid),
    .io_to_pes_25_out_bits(PENetwork_18_io_to_pes_25_out_bits),
    .io_to_pes_26_in_valid(PENetwork_18_io_to_pes_26_in_valid),
    .io_to_pes_26_in_bits(PENetwork_18_io_to_pes_26_in_bits),
    .io_to_pes_26_out_valid(PENetwork_18_io_to_pes_26_out_valid),
    .io_to_pes_26_out_bits(PENetwork_18_io_to_pes_26_out_bits),
    .io_to_pes_27_in_valid(PENetwork_18_io_to_pes_27_in_valid),
    .io_to_pes_27_in_bits(PENetwork_18_io_to_pes_27_in_bits),
    .io_to_pes_27_out_valid(PENetwork_18_io_to_pes_27_out_valid),
    .io_to_pes_27_out_bits(PENetwork_18_io_to_pes_27_out_bits),
    .io_to_pes_28_in_valid(PENetwork_18_io_to_pes_28_in_valid),
    .io_to_pes_28_in_bits(PENetwork_18_io_to_pes_28_in_bits),
    .io_to_pes_28_out_valid(PENetwork_18_io_to_pes_28_out_valid),
    .io_to_pes_28_out_bits(PENetwork_18_io_to_pes_28_out_bits),
    .io_to_pes_29_in_valid(PENetwork_18_io_to_pes_29_in_valid),
    .io_to_pes_29_in_bits(PENetwork_18_io_to_pes_29_in_bits),
    .io_to_mem_valid(PENetwork_18_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_18_io_to_mem_bits)
  );
  PENetwork PENetwork_19 ( // @[pe.scala 229:13]
    .io_to_pes_0_in_valid(PENetwork_19_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_19_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_19_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_19_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_19_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_19_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_19_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_19_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_19_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_19_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_19_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_19_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_19_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_19_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_19_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_19_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_19_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_19_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_19_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_19_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_19_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_19_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_19_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_19_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_19_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_19_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_19_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_19_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_19_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_19_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_19_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_19_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_19_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_19_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_19_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_19_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_19_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_19_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_19_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_19_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_19_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_19_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_19_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_19_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_19_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_19_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_19_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_19_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_19_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_19_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_19_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_19_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_19_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_19_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_19_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_19_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_19_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_19_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_19_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_19_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_19_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_19_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_19_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_19_io_to_pes_15_out_bits),
    .io_to_pes_16_in_valid(PENetwork_19_io_to_pes_16_in_valid),
    .io_to_pes_16_in_bits(PENetwork_19_io_to_pes_16_in_bits),
    .io_to_pes_16_out_valid(PENetwork_19_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_19_io_to_pes_16_out_bits),
    .io_to_pes_17_in_valid(PENetwork_19_io_to_pes_17_in_valid),
    .io_to_pes_17_in_bits(PENetwork_19_io_to_pes_17_in_bits),
    .io_to_pes_17_out_valid(PENetwork_19_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_19_io_to_pes_17_out_bits),
    .io_to_pes_18_in_valid(PENetwork_19_io_to_pes_18_in_valid),
    .io_to_pes_18_in_bits(PENetwork_19_io_to_pes_18_in_bits),
    .io_to_pes_18_out_valid(PENetwork_19_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_19_io_to_pes_18_out_bits),
    .io_to_pes_19_in_valid(PENetwork_19_io_to_pes_19_in_valid),
    .io_to_pes_19_in_bits(PENetwork_19_io_to_pes_19_in_bits),
    .io_to_pes_19_out_valid(PENetwork_19_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_19_io_to_pes_19_out_bits),
    .io_to_pes_20_in_valid(PENetwork_19_io_to_pes_20_in_valid),
    .io_to_pes_20_in_bits(PENetwork_19_io_to_pes_20_in_bits),
    .io_to_pes_20_out_valid(PENetwork_19_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_19_io_to_pes_20_out_bits),
    .io_to_pes_21_in_valid(PENetwork_19_io_to_pes_21_in_valid),
    .io_to_pes_21_in_bits(PENetwork_19_io_to_pes_21_in_bits),
    .io_to_pes_21_out_valid(PENetwork_19_io_to_pes_21_out_valid),
    .io_to_pes_21_out_bits(PENetwork_19_io_to_pes_21_out_bits),
    .io_to_pes_22_in_valid(PENetwork_19_io_to_pes_22_in_valid),
    .io_to_pes_22_in_bits(PENetwork_19_io_to_pes_22_in_bits),
    .io_to_pes_22_out_valid(PENetwork_19_io_to_pes_22_out_valid),
    .io_to_pes_22_out_bits(PENetwork_19_io_to_pes_22_out_bits),
    .io_to_pes_23_in_valid(PENetwork_19_io_to_pes_23_in_valid),
    .io_to_pes_23_in_bits(PENetwork_19_io_to_pes_23_in_bits),
    .io_to_pes_23_out_valid(PENetwork_19_io_to_pes_23_out_valid),
    .io_to_pes_23_out_bits(PENetwork_19_io_to_pes_23_out_bits),
    .io_to_pes_24_in_valid(PENetwork_19_io_to_pes_24_in_valid),
    .io_to_pes_24_in_bits(PENetwork_19_io_to_pes_24_in_bits),
    .io_to_pes_24_out_valid(PENetwork_19_io_to_pes_24_out_valid),
    .io_to_pes_24_out_bits(PENetwork_19_io_to_pes_24_out_bits),
    .io_to_pes_25_in_valid(PENetwork_19_io_to_pes_25_in_valid),
    .io_to_pes_25_in_bits(PENetwork_19_io_to_pes_25_in_bits),
    .io_to_pes_25_out_valid(PENetwork_19_io_to_pes_25_out_valid),
    .io_to_pes_25_out_bits(PENetwork_19_io_to_pes_25_out_bits),
    .io_to_pes_26_in_valid(PENetwork_19_io_to_pes_26_in_valid),
    .io_to_pes_26_in_bits(PENetwork_19_io_to_pes_26_in_bits),
    .io_to_pes_26_out_valid(PENetwork_19_io_to_pes_26_out_valid),
    .io_to_pes_26_out_bits(PENetwork_19_io_to_pes_26_out_bits),
    .io_to_pes_27_in_valid(PENetwork_19_io_to_pes_27_in_valid),
    .io_to_pes_27_in_bits(PENetwork_19_io_to_pes_27_in_bits),
    .io_to_pes_27_out_valid(PENetwork_19_io_to_pes_27_out_valid),
    .io_to_pes_27_out_bits(PENetwork_19_io_to_pes_27_out_bits),
    .io_to_pes_28_in_valid(PENetwork_19_io_to_pes_28_in_valid),
    .io_to_pes_28_in_bits(PENetwork_19_io_to_pes_28_in_bits),
    .io_to_pes_28_out_valid(PENetwork_19_io_to_pes_28_out_valid),
    .io_to_pes_28_out_bits(PENetwork_19_io_to_pes_28_out_bits),
    .io_to_pes_29_in_valid(PENetwork_19_io_to_pes_29_in_valid),
    .io_to_pes_29_in_bits(PENetwork_19_io_to_pes_29_in_bits),
    .io_to_mem_valid(PENetwork_19_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_19_io_to_mem_bits)
  );
  PENetwork PENetwork_20 ( // @[pe.scala 229:13]
    .io_to_pes_0_in_valid(PENetwork_20_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_20_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_20_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_20_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_20_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_20_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_20_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_20_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_20_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_20_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_20_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_20_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_20_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_20_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_20_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_20_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_20_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_20_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_20_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_20_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_20_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_20_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_20_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_20_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_20_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_20_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_20_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_20_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_20_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_20_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_20_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_20_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_20_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_20_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_20_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_20_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_20_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_20_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_20_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_20_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_20_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_20_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_20_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_20_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_20_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_20_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_20_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_20_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_20_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_20_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_20_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_20_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_20_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_20_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_20_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_20_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_20_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_20_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_20_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_20_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_20_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_20_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_20_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_20_io_to_pes_15_out_bits),
    .io_to_pes_16_in_valid(PENetwork_20_io_to_pes_16_in_valid),
    .io_to_pes_16_in_bits(PENetwork_20_io_to_pes_16_in_bits),
    .io_to_pes_16_out_valid(PENetwork_20_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_20_io_to_pes_16_out_bits),
    .io_to_pes_17_in_valid(PENetwork_20_io_to_pes_17_in_valid),
    .io_to_pes_17_in_bits(PENetwork_20_io_to_pes_17_in_bits),
    .io_to_pes_17_out_valid(PENetwork_20_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_20_io_to_pes_17_out_bits),
    .io_to_pes_18_in_valid(PENetwork_20_io_to_pes_18_in_valid),
    .io_to_pes_18_in_bits(PENetwork_20_io_to_pes_18_in_bits),
    .io_to_pes_18_out_valid(PENetwork_20_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_20_io_to_pes_18_out_bits),
    .io_to_pes_19_in_valid(PENetwork_20_io_to_pes_19_in_valid),
    .io_to_pes_19_in_bits(PENetwork_20_io_to_pes_19_in_bits),
    .io_to_pes_19_out_valid(PENetwork_20_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_20_io_to_pes_19_out_bits),
    .io_to_pes_20_in_valid(PENetwork_20_io_to_pes_20_in_valid),
    .io_to_pes_20_in_bits(PENetwork_20_io_to_pes_20_in_bits),
    .io_to_pes_20_out_valid(PENetwork_20_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_20_io_to_pes_20_out_bits),
    .io_to_pes_21_in_valid(PENetwork_20_io_to_pes_21_in_valid),
    .io_to_pes_21_in_bits(PENetwork_20_io_to_pes_21_in_bits),
    .io_to_pes_21_out_valid(PENetwork_20_io_to_pes_21_out_valid),
    .io_to_pes_21_out_bits(PENetwork_20_io_to_pes_21_out_bits),
    .io_to_pes_22_in_valid(PENetwork_20_io_to_pes_22_in_valid),
    .io_to_pes_22_in_bits(PENetwork_20_io_to_pes_22_in_bits),
    .io_to_pes_22_out_valid(PENetwork_20_io_to_pes_22_out_valid),
    .io_to_pes_22_out_bits(PENetwork_20_io_to_pes_22_out_bits),
    .io_to_pes_23_in_valid(PENetwork_20_io_to_pes_23_in_valid),
    .io_to_pes_23_in_bits(PENetwork_20_io_to_pes_23_in_bits),
    .io_to_pes_23_out_valid(PENetwork_20_io_to_pes_23_out_valid),
    .io_to_pes_23_out_bits(PENetwork_20_io_to_pes_23_out_bits),
    .io_to_pes_24_in_valid(PENetwork_20_io_to_pes_24_in_valid),
    .io_to_pes_24_in_bits(PENetwork_20_io_to_pes_24_in_bits),
    .io_to_pes_24_out_valid(PENetwork_20_io_to_pes_24_out_valid),
    .io_to_pes_24_out_bits(PENetwork_20_io_to_pes_24_out_bits),
    .io_to_pes_25_in_valid(PENetwork_20_io_to_pes_25_in_valid),
    .io_to_pes_25_in_bits(PENetwork_20_io_to_pes_25_in_bits),
    .io_to_pes_25_out_valid(PENetwork_20_io_to_pes_25_out_valid),
    .io_to_pes_25_out_bits(PENetwork_20_io_to_pes_25_out_bits),
    .io_to_pes_26_in_valid(PENetwork_20_io_to_pes_26_in_valid),
    .io_to_pes_26_in_bits(PENetwork_20_io_to_pes_26_in_bits),
    .io_to_pes_26_out_valid(PENetwork_20_io_to_pes_26_out_valid),
    .io_to_pes_26_out_bits(PENetwork_20_io_to_pes_26_out_bits),
    .io_to_pes_27_in_valid(PENetwork_20_io_to_pes_27_in_valid),
    .io_to_pes_27_in_bits(PENetwork_20_io_to_pes_27_in_bits),
    .io_to_pes_27_out_valid(PENetwork_20_io_to_pes_27_out_valid),
    .io_to_pes_27_out_bits(PENetwork_20_io_to_pes_27_out_bits),
    .io_to_pes_28_in_valid(PENetwork_20_io_to_pes_28_in_valid),
    .io_to_pes_28_in_bits(PENetwork_20_io_to_pes_28_in_bits),
    .io_to_pes_28_out_valid(PENetwork_20_io_to_pes_28_out_valid),
    .io_to_pes_28_out_bits(PENetwork_20_io_to_pes_28_out_bits),
    .io_to_pes_29_in_valid(PENetwork_20_io_to_pes_29_in_valid),
    .io_to_pes_29_in_bits(PENetwork_20_io_to_pes_29_in_bits),
    .io_to_mem_valid(PENetwork_20_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_20_io_to_mem_bits)
  );
  PENetwork PENetwork_21 ( // @[pe.scala 229:13]
    .io_to_pes_0_in_valid(PENetwork_21_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_21_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_21_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_21_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_21_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_21_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_21_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_21_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_21_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_21_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_21_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_21_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_21_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_21_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_21_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_21_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_21_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_21_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_21_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_21_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_21_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_21_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_21_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_21_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_21_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_21_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_21_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_21_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_21_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_21_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_21_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_21_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_21_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_21_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_21_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_21_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_21_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_21_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_21_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_21_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_21_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_21_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_21_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_21_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_21_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_21_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_21_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_21_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_21_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_21_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_21_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_21_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_21_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_21_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_21_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_21_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_21_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_21_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_21_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_21_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_21_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_21_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_21_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_21_io_to_pes_15_out_bits),
    .io_to_pes_16_in_valid(PENetwork_21_io_to_pes_16_in_valid),
    .io_to_pes_16_in_bits(PENetwork_21_io_to_pes_16_in_bits),
    .io_to_pes_16_out_valid(PENetwork_21_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_21_io_to_pes_16_out_bits),
    .io_to_pes_17_in_valid(PENetwork_21_io_to_pes_17_in_valid),
    .io_to_pes_17_in_bits(PENetwork_21_io_to_pes_17_in_bits),
    .io_to_pes_17_out_valid(PENetwork_21_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_21_io_to_pes_17_out_bits),
    .io_to_pes_18_in_valid(PENetwork_21_io_to_pes_18_in_valid),
    .io_to_pes_18_in_bits(PENetwork_21_io_to_pes_18_in_bits),
    .io_to_pes_18_out_valid(PENetwork_21_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_21_io_to_pes_18_out_bits),
    .io_to_pes_19_in_valid(PENetwork_21_io_to_pes_19_in_valid),
    .io_to_pes_19_in_bits(PENetwork_21_io_to_pes_19_in_bits),
    .io_to_pes_19_out_valid(PENetwork_21_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_21_io_to_pes_19_out_bits),
    .io_to_pes_20_in_valid(PENetwork_21_io_to_pes_20_in_valid),
    .io_to_pes_20_in_bits(PENetwork_21_io_to_pes_20_in_bits),
    .io_to_pes_20_out_valid(PENetwork_21_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_21_io_to_pes_20_out_bits),
    .io_to_pes_21_in_valid(PENetwork_21_io_to_pes_21_in_valid),
    .io_to_pes_21_in_bits(PENetwork_21_io_to_pes_21_in_bits),
    .io_to_pes_21_out_valid(PENetwork_21_io_to_pes_21_out_valid),
    .io_to_pes_21_out_bits(PENetwork_21_io_to_pes_21_out_bits),
    .io_to_pes_22_in_valid(PENetwork_21_io_to_pes_22_in_valid),
    .io_to_pes_22_in_bits(PENetwork_21_io_to_pes_22_in_bits),
    .io_to_pes_22_out_valid(PENetwork_21_io_to_pes_22_out_valid),
    .io_to_pes_22_out_bits(PENetwork_21_io_to_pes_22_out_bits),
    .io_to_pes_23_in_valid(PENetwork_21_io_to_pes_23_in_valid),
    .io_to_pes_23_in_bits(PENetwork_21_io_to_pes_23_in_bits),
    .io_to_pes_23_out_valid(PENetwork_21_io_to_pes_23_out_valid),
    .io_to_pes_23_out_bits(PENetwork_21_io_to_pes_23_out_bits),
    .io_to_pes_24_in_valid(PENetwork_21_io_to_pes_24_in_valid),
    .io_to_pes_24_in_bits(PENetwork_21_io_to_pes_24_in_bits),
    .io_to_pes_24_out_valid(PENetwork_21_io_to_pes_24_out_valid),
    .io_to_pes_24_out_bits(PENetwork_21_io_to_pes_24_out_bits),
    .io_to_pes_25_in_valid(PENetwork_21_io_to_pes_25_in_valid),
    .io_to_pes_25_in_bits(PENetwork_21_io_to_pes_25_in_bits),
    .io_to_pes_25_out_valid(PENetwork_21_io_to_pes_25_out_valid),
    .io_to_pes_25_out_bits(PENetwork_21_io_to_pes_25_out_bits),
    .io_to_pes_26_in_valid(PENetwork_21_io_to_pes_26_in_valid),
    .io_to_pes_26_in_bits(PENetwork_21_io_to_pes_26_in_bits),
    .io_to_pes_26_out_valid(PENetwork_21_io_to_pes_26_out_valid),
    .io_to_pes_26_out_bits(PENetwork_21_io_to_pes_26_out_bits),
    .io_to_pes_27_in_valid(PENetwork_21_io_to_pes_27_in_valid),
    .io_to_pes_27_in_bits(PENetwork_21_io_to_pes_27_in_bits),
    .io_to_pes_27_out_valid(PENetwork_21_io_to_pes_27_out_valid),
    .io_to_pes_27_out_bits(PENetwork_21_io_to_pes_27_out_bits),
    .io_to_pes_28_in_valid(PENetwork_21_io_to_pes_28_in_valid),
    .io_to_pes_28_in_bits(PENetwork_21_io_to_pes_28_in_bits),
    .io_to_pes_28_out_valid(PENetwork_21_io_to_pes_28_out_valid),
    .io_to_pes_28_out_bits(PENetwork_21_io_to_pes_28_out_bits),
    .io_to_pes_29_in_valid(PENetwork_21_io_to_pes_29_in_valid),
    .io_to_pes_29_in_bits(PENetwork_21_io_to_pes_29_in_bits),
    .io_to_mem_valid(PENetwork_21_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_21_io_to_mem_bits)
  );
  PENetwork_22 PENetwork_22 ( // @[pe.scala 229:13]
    .io_to_pes_0_in_valid(PENetwork_22_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_22_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_22_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_22_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_22_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_22_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_22_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_22_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_22_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_22_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_22_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_22_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_22_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_22_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_22_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_22_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_22_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_22_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_22_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_22_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_22_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_22_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_22_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_22_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_22_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_22_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_22_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_22_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_22_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_22_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_22_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_22_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_22_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_22_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_22_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_22_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_22_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_22_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_22_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_22_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_22_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_22_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_22_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_22_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_22_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_22_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_22_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_22_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_22_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_22_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_22_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_22_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_22_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_22_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_22_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_22_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_22_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_22_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_22_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_22_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_22_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_22_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_22_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_22_io_to_pes_15_out_bits),
    .io_to_pes_16_in_valid(PENetwork_22_io_to_pes_16_in_valid),
    .io_to_pes_16_in_bits(PENetwork_22_io_to_pes_16_in_bits),
    .io_to_pes_16_out_valid(PENetwork_22_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_22_io_to_pes_16_out_bits),
    .io_to_pes_17_in_valid(PENetwork_22_io_to_pes_17_in_valid),
    .io_to_pes_17_in_bits(PENetwork_22_io_to_pes_17_in_bits),
    .io_to_pes_17_out_valid(PENetwork_22_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_22_io_to_pes_17_out_bits),
    .io_to_pes_18_in_valid(PENetwork_22_io_to_pes_18_in_valid),
    .io_to_pes_18_in_bits(PENetwork_22_io_to_pes_18_in_bits),
    .io_to_pes_18_out_valid(PENetwork_22_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_22_io_to_pes_18_out_bits),
    .io_to_pes_19_in_valid(PENetwork_22_io_to_pes_19_in_valid),
    .io_to_pes_19_in_bits(PENetwork_22_io_to_pes_19_in_bits),
    .io_to_pes_19_out_valid(PENetwork_22_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_22_io_to_pes_19_out_bits),
    .io_to_pes_20_in_valid(PENetwork_22_io_to_pes_20_in_valid),
    .io_to_pes_20_in_bits(PENetwork_22_io_to_pes_20_in_bits),
    .io_to_pes_20_out_valid(PENetwork_22_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_22_io_to_pes_20_out_bits),
    .io_to_pes_21_in_valid(PENetwork_22_io_to_pes_21_in_valid),
    .io_to_pes_21_in_bits(PENetwork_22_io_to_pes_21_in_bits),
    .io_to_mem_valid(PENetwork_22_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_22_io_to_mem_bits)
  );
  PENetwork_22 PENetwork_23 ( // @[pe.scala 229:13]
    .io_to_pes_0_in_valid(PENetwork_23_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_23_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_23_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_23_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_23_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_23_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_23_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_23_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_23_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_23_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_23_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_23_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_23_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_23_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_23_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_23_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_23_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_23_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_23_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_23_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_23_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_23_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_23_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_23_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_23_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_23_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_23_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_23_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_23_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_23_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_23_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_23_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_23_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_23_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_23_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_23_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_23_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_23_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_23_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_23_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_23_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_23_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_23_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_23_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_23_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_23_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_23_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_23_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_23_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_23_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_23_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_23_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_23_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_23_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_23_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_23_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_23_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_23_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_23_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_23_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_23_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_23_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_23_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_23_io_to_pes_15_out_bits),
    .io_to_pes_16_in_valid(PENetwork_23_io_to_pes_16_in_valid),
    .io_to_pes_16_in_bits(PENetwork_23_io_to_pes_16_in_bits),
    .io_to_pes_16_out_valid(PENetwork_23_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_23_io_to_pes_16_out_bits),
    .io_to_pes_17_in_valid(PENetwork_23_io_to_pes_17_in_valid),
    .io_to_pes_17_in_bits(PENetwork_23_io_to_pes_17_in_bits),
    .io_to_pes_17_out_valid(PENetwork_23_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_23_io_to_pes_17_out_bits),
    .io_to_pes_18_in_valid(PENetwork_23_io_to_pes_18_in_valid),
    .io_to_pes_18_in_bits(PENetwork_23_io_to_pes_18_in_bits),
    .io_to_pes_18_out_valid(PENetwork_23_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_23_io_to_pes_18_out_bits),
    .io_to_pes_19_in_valid(PENetwork_23_io_to_pes_19_in_valid),
    .io_to_pes_19_in_bits(PENetwork_23_io_to_pes_19_in_bits),
    .io_to_pes_19_out_valid(PENetwork_23_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_23_io_to_pes_19_out_bits),
    .io_to_pes_20_in_valid(PENetwork_23_io_to_pes_20_in_valid),
    .io_to_pes_20_in_bits(PENetwork_23_io_to_pes_20_in_bits),
    .io_to_pes_20_out_valid(PENetwork_23_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_23_io_to_pes_20_out_bits),
    .io_to_pes_21_in_valid(PENetwork_23_io_to_pes_21_in_valid),
    .io_to_pes_21_in_bits(PENetwork_23_io_to_pes_21_in_bits),
    .io_to_mem_valid(PENetwork_23_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_23_io_to_mem_bits)
  );
  PENetwork_22 PENetwork_24 ( // @[pe.scala 229:13]
    .io_to_pes_0_in_valid(PENetwork_24_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_24_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_24_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_24_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_24_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_24_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_24_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_24_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_24_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_24_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_24_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_24_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_24_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_24_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_24_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_24_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_24_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_24_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_24_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_24_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_24_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_24_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_24_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_24_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_24_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_24_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_24_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_24_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_24_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_24_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_24_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_24_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_24_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_24_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_24_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_24_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_24_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_24_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_24_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_24_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_24_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_24_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_24_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_24_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_24_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_24_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_24_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_24_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_24_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_24_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_24_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_24_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_24_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_24_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_24_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_24_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_24_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_24_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_24_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_24_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_24_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_24_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_24_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_24_io_to_pes_15_out_bits),
    .io_to_pes_16_in_valid(PENetwork_24_io_to_pes_16_in_valid),
    .io_to_pes_16_in_bits(PENetwork_24_io_to_pes_16_in_bits),
    .io_to_pes_16_out_valid(PENetwork_24_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_24_io_to_pes_16_out_bits),
    .io_to_pes_17_in_valid(PENetwork_24_io_to_pes_17_in_valid),
    .io_to_pes_17_in_bits(PENetwork_24_io_to_pes_17_in_bits),
    .io_to_pes_17_out_valid(PENetwork_24_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_24_io_to_pes_17_out_bits),
    .io_to_pes_18_in_valid(PENetwork_24_io_to_pes_18_in_valid),
    .io_to_pes_18_in_bits(PENetwork_24_io_to_pes_18_in_bits),
    .io_to_pes_18_out_valid(PENetwork_24_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_24_io_to_pes_18_out_bits),
    .io_to_pes_19_in_valid(PENetwork_24_io_to_pes_19_in_valid),
    .io_to_pes_19_in_bits(PENetwork_24_io_to_pes_19_in_bits),
    .io_to_pes_19_out_valid(PENetwork_24_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_24_io_to_pes_19_out_bits),
    .io_to_pes_20_in_valid(PENetwork_24_io_to_pes_20_in_valid),
    .io_to_pes_20_in_bits(PENetwork_24_io_to_pes_20_in_bits),
    .io_to_pes_20_out_valid(PENetwork_24_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_24_io_to_pes_20_out_bits),
    .io_to_pes_21_in_valid(PENetwork_24_io_to_pes_21_in_valid),
    .io_to_pes_21_in_bits(PENetwork_24_io_to_pes_21_in_bits),
    .io_to_mem_valid(PENetwork_24_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_24_io_to_mem_bits)
  );
  PENetwork_22 PENetwork_25 ( // @[pe.scala 229:13]
    .io_to_pes_0_in_valid(PENetwork_25_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_25_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_25_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_25_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_25_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_25_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_25_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_25_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_25_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_25_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_25_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_25_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_25_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_25_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_25_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_25_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_25_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_25_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_25_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_25_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_25_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_25_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_25_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_25_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_25_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_25_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_25_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_25_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_25_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_25_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_25_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_25_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_25_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_25_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_25_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_25_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_25_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_25_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_25_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_25_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_25_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_25_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_25_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_25_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_25_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_25_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_25_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_25_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_25_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_25_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_25_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_25_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_25_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_25_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_25_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_25_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_25_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_25_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_25_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_25_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_25_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_25_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_25_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_25_io_to_pes_15_out_bits),
    .io_to_pes_16_in_valid(PENetwork_25_io_to_pes_16_in_valid),
    .io_to_pes_16_in_bits(PENetwork_25_io_to_pes_16_in_bits),
    .io_to_pes_16_out_valid(PENetwork_25_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_25_io_to_pes_16_out_bits),
    .io_to_pes_17_in_valid(PENetwork_25_io_to_pes_17_in_valid),
    .io_to_pes_17_in_bits(PENetwork_25_io_to_pes_17_in_bits),
    .io_to_pes_17_out_valid(PENetwork_25_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_25_io_to_pes_17_out_bits),
    .io_to_pes_18_in_valid(PENetwork_25_io_to_pes_18_in_valid),
    .io_to_pes_18_in_bits(PENetwork_25_io_to_pes_18_in_bits),
    .io_to_pes_18_out_valid(PENetwork_25_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_25_io_to_pes_18_out_bits),
    .io_to_pes_19_in_valid(PENetwork_25_io_to_pes_19_in_valid),
    .io_to_pes_19_in_bits(PENetwork_25_io_to_pes_19_in_bits),
    .io_to_pes_19_out_valid(PENetwork_25_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_25_io_to_pes_19_out_bits),
    .io_to_pes_20_in_valid(PENetwork_25_io_to_pes_20_in_valid),
    .io_to_pes_20_in_bits(PENetwork_25_io_to_pes_20_in_bits),
    .io_to_pes_20_out_valid(PENetwork_25_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_25_io_to_pes_20_out_bits),
    .io_to_pes_21_in_valid(PENetwork_25_io_to_pes_21_in_valid),
    .io_to_pes_21_in_bits(PENetwork_25_io_to_pes_21_in_bits),
    .io_to_mem_valid(PENetwork_25_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_25_io_to_mem_bits)
  );
  PENetwork_22 PENetwork_26 ( // @[pe.scala 229:13]
    .io_to_pes_0_in_valid(PENetwork_26_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_26_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_26_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_26_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_26_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_26_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_26_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_26_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_26_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_26_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_26_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_26_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_26_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_26_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_26_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_26_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_26_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_26_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_26_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_26_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_26_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_26_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_26_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_26_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_26_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_26_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_26_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_26_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_26_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_26_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_26_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_26_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_26_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_26_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_26_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_26_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_26_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_26_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_26_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_26_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_26_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_26_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_26_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_26_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_26_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_26_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_26_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_26_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_26_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_26_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_26_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_26_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_26_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_26_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_26_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_26_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_26_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_26_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_26_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_26_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_26_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_26_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_26_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_26_io_to_pes_15_out_bits),
    .io_to_pes_16_in_valid(PENetwork_26_io_to_pes_16_in_valid),
    .io_to_pes_16_in_bits(PENetwork_26_io_to_pes_16_in_bits),
    .io_to_pes_16_out_valid(PENetwork_26_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_26_io_to_pes_16_out_bits),
    .io_to_pes_17_in_valid(PENetwork_26_io_to_pes_17_in_valid),
    .io_to_pes_17_in_bits(PENetwork_26_io_to_pes_17_in_bits),
    .io_to_pes_17_out_valid(PENetwork_26_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_26_io_to_pes_17_out_bits),
    .io_to_pes_18_in_valid(PENetwork_26_io_to_pes_18_in_valid),
    .io_to_pes_18_in_bits(PENetwork_26_io_to_pes_18_in_bits),
    .io_to_pes_18_out_valid(PENetwork_26_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_26_io_to_pes_18_out_bits),
    .io_to_pes_19_in_valid(PENetwork_26_io_to_pes_19_in_valid),
    .io_to_pes_19_in_bits(PENetwork_26_io_to_pes_19_in_bits),
    .io_to_pes_19_out_valid(PENetwork_26_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_26_io_to_pes_19_out_bits),
    .io_to_pes_20_in_valid(PENetwork_26_io_to_pes_20_in_valid),
    .io_to_pes_20_in_bits(PENetwork_26_io_to_pes_20_in_bits),
    .io_to_pes_20_out_valid(PENetwork_26_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_26_io_to_pes_20_out_bits),
    .io_to_pes_21_in_valid(PENetwork_26_io_to_pes_21_in_valid),
    .io_to_pes_21_in_bits(PENetwork_26_io_to_pes_21_in_bits),
    .io_to_mem_valid(PENetwork_26_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_26_io_to_mem_bits)
  );
  PENetwork_22 PENetwork_27 ( // @[pe.scala 229:13]
    .io_to_pes_0_in_valid(PENetwork_27_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_27_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_27_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_27_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_27_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_27_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_27_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_27_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_27_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_27_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_27_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_27_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_27_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_27_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_27_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_27_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_27_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_27_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_27_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_27_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_27_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_27_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_27_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_27_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_27_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_27_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_27_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_27_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_27_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_27_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_27_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_27_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_27_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_27_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_27_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_27_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_27_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_27_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_27_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_27_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_27_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_27_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_27_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_27_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_27_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_27_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_27_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_27_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_27_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_27_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_27_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_27_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_27_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_27_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_27_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_27_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_27_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_27_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_27_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_27_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_27_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_27_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_27_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_27_io_to_pes_15_out_bits),
    .io_to_pes_16_in_valid(PENetwork_27_io_to_pes_16_in_valid),
    .io_to_pes_16_in_bits(PENetwork_27_io_to_pes_16_in_bits),
    .io_to_pes_16_out_valid(PENetwork_27_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_27_io_to_pes_16_out_bits),
    .io_to_pes_17_in_valid(PENetwork_27_io_to_pes_17_in_valid),
    .io_to_pes_17_in_bits(PENetwork_27_io_to_pes_17_in_bits),
    .io_to_pes_17_out_valid(PENetwork_27_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_27_io_to_pes_17_out_bits),
    .io_to_pes_18_in_valid(PENetwork_27_io_to_pes_18_in_valid),
    .io_to_pes_18_in_bits(PENetwork_27_io_to_pes_18_in_bits),
    .io_to_pes_18_out_valid(PENetwork_27_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_27_io_to_pes_18_out_bits),
    .io_to_pes_19_in_valid(PENetwork_27_io_to_pes_19_in_valid),
    .io_to_pes_19_in_bits(PENetwork_27_io_to_pes_19_in_bits),
    .io_to_pes_19_out_valid(PENetwork_27_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_27_io_to_pes_19_out_bits),
    .io_to_pes_20_in_valid(PENetwork_27_io_to_pes_20_in_valid),
    .io_to_pes_20_in_bits(PENetwork_27_io_to_pes_20_in_bits),
    .io_to_pes_20_out_valid(PENetwork_27_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_27_io_to_pes_20_out_bits),
    .io_to_pes_21_in_valid(PENetwork_27_io_to_pes_21_in_valid),
    .io_to_pes_21_in_bits(PENetwork_27_io_to_pes_21_in_bits),
    .io_to_mem_valid(PENetwork_27_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_27_io_to_mem_bits)
  );
  PENetwork_22 PENetwork_28 ( // @[pe.scala 229:13]
    .io_to_pes_0_in_valid(PENetwork_28_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_28_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_28_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_28_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_28_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_28_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_28_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_28_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_28_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_28_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_28_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_28_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_28_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_28_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_28_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_28_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_28_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_28_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_28_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_28_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_28_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_28_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_28_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_28_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_28_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_28_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_28_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_28_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_28_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_28_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_28_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_28_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_28_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_28_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_28_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_28_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_28_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_28_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_28_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_28_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_28_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_28_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_28_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_28_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_28_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_28_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_28_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_28_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_28_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_28_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_28_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_28_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_28_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_28_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_28_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_28_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_28_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_28_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_28_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_28_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_28_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_28_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_28_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_28_io_to_pes_15_out_bits),
    .io_to_pes_16_in_valid(PENetwork_28_io_to_pes_16_in_valid),
    .io_to_pes_16_in_bits(PENetwork_28_io_to_pes_16_in_bits),
    .io_to_pes_16_out_valid(PENetwork_28_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_28_io_to_pes_16_out_bits),
    .io_to_pes_17_in_valid(PENetwork_28_io_to_pes_17_in_valid),
    .io_to_pes_17_in_bits(PENetwork_28_io_to_pes_17_in_bits),
    .io_to_pes_17_out_valid(PENetwork_28_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_28_io_to_pes_17_out_bits),
    .io_to_pes_18_in_valid(PENetwork_28_io_to_pes_18_in_valid),
    .io_to_pes_18_in_bits(PENetwork_28_io_to_pes_18_in_bits),
    .io_to_pes_18_out_valid(PENetwork_28_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_28_io_to_pes_18_out_bits),
    .io_to_pes_19_in_valid(PENetwork_28_io_to_pes_19_in_valid),
    .io_to_pes_19_in_bits(PENetwork_28_io_to_pes_19_in_bits),
    .io_to_pes_19_out_valid(PENetwork_28_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_28_io_to_pes_19_out_bits),
    .io_to_pes_20_in_valid(PENetwork_28_io_to_pes_20_in_valid),
    .io_to_pes_20_in_bits(PENetwork_28_io_to_pes_20_in_bits),
    .io_to_pes_20_out_valid(PENetwork_28_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_28_io_to_pes_20_out_bits),
    .io_to_pes_21_in_valid(PENetwork_28_io_to_pes_21_in_valid),
    .io_to_pes_21_in_bits(PENetwork_28_io_to_pes_21_in_bits),
    .io_to_mem_valid(PENetwork_28_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_28_io_to_mem_bits)
  );
  PENetwork_22 PENetwork_29 ( // @[pe.scala 229:13]
    .io_to_pes_0_in_valid(PENetwork_29_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_29_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_29_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_29_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_29_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_29_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_29_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_29_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_29_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_29_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_29_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_29_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_29_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_29_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_29_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_29_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_29_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_29_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_29_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_29_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_29_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_29_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_29_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_29_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_29_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_29_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_29_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_29_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_29_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_29_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_29_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_29_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_29_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_29_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_29_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_29_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_29_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_29_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_29_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_29_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_29_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_29_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_29_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_29_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_29_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_29_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_29_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_29_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_29_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_29_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_29_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_29_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_29_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_29_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_29_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_29_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_29_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_29_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_29_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_29_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_29_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_29_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_29_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_29_io_to_pes_15_out_bits),
    .io_to_pes_16_in_valid(PENetwork_29_io_to_pes_16_in_valid),
    .io_to_pes_16_in_bits(PENetwork_29_io_to_pes_16_in_bits),
    .io_to_pes_16_out_valid(PENetwork_29_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_29_io_to_pes_16_out_bits),
    .io_to_pes_17_in_valid(PENetwork_29_io_to_pes_17_in_valid),
    .io_to_pes_17_in_bits(PENetwork_29_io_to_pes_17_in_bits),
    .io_to_pes_17_out_valid(PENetwork_29_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_29_io_to_pes_17_out_bits),
    .io_to_pes_18_in_valid(PENetwork_29_io_to_pes_18_in_valid),
    .io_to_pes_18_in_bits(PENetwork_29_io_to_pes_18_in_bits),
    .io_to_pes_18_out_valid(PENetwork_29_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_29_io_to_pes_18_out_bits),
    .io_to_pes_19_in_valid(PENetwork_29_io_to_pes_19_in_valid),
    .io_to_pes_19_in_bits(PENetwork_29_io_to_pes_19_in_bits),
    .io_to_pes_19_out_valid(PENetwork_29_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_29_io_to_pes_19_out_bits),
    .io_to_pes_20_in_valid(PENetwork_29_io_to_pes_20_in_valid),
    .io_to_pes_20_in_bits(PENetwork_29_io_to_pes_20_in_bits),
    .io_to_pes_20_out_valid(PENetwork_29_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_29_io_to_pes_20_out_bits),
    .io_to_pes_21_in_valid(PENetwork_29_io_to_pes_21_in_valid),
    .io_to_pes_21_in_bits(PENetwork_29_io_to_pes_21_in_bits),
    .io_to_mem_valid(PENetwork_29_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_29_io_to_mem_bits)
  );
  PENetwork_22 PENetwork_30 ( // @[pe.scala 229:13]
    .io_to_pes_0_in_valid(PENetwork_30_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_30_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_30_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_30_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_30_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_30_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_30_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_30_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_30_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_30_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_30_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_30_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_30_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_30_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_30_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_30_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_30_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_30_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_30_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_30_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_30_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_30_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_30_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_30_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_30_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_30_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_30_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_30_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_30_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_30_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_30_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_30_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_30_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_30_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_30_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_30_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_30_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_30_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_30_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_30_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_30_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_30_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_30_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_30_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_30_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_30_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_30_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_30_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_30_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_30_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_30_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_30_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_30_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_30_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_30_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_30_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_30_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_30_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_30_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_30_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_30_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_30_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_30_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_30_io_to_pes_15_out_bits),
    .io_to_pes_16_in_valid(PENetwork_30_io_to_pes_16_in_valid),
    .io_to_pes_16_in_bits(PENetwork_30_io_to_pes_16_in_bits),
    .io_to_pes_16_out_valid(PENetwork_30_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_30_io_to_pes_16_out_bits),
    .io_to_pes_17_in_valid(PENetwork_30_io_to_pes_17_in_valid),
    .io_to_pes_17_in_bits(PENetwork_30_io_to_pes_17_in_bits),
    .io_to_pes_17_out_valid(PENetwork_30_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_30_io_to_pes_17_out_bits),
    .io_to_pes_18_in_valid(PENetwork_30_io_to_pes_18_in_valid),
    .io_to_pes_18_in_bits(PENetwork_30_io_to_pes_18_in_bits),
    .io_to_pes_18_out_valid(PENetwork_30_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_30_io_to_pes_18_out_bits),
    .io_to_pes_19_in_valid(PENetwork_30_io_to_pes_19_in_valid),
    .io_to_pes_19_in_bits(PENetwork_30_io_to_pes_19_in_bits),
    .io_to_pes_19_out_valid(PENetwork_30_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_30_io_to_pes_19_out_bits),
    .io_to_pes_20_in_valid(PENetwork_30_io_to_pes_20_in_valid),
    .io_to_pes_20_in_bits(PENetwork_30_io_to_pes_20_in_bits),
    .io_to_pes_20_out_valid(PENetwork_30_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_30_io_to_pes_20_out_bits),
    .io_to_pes_21_in_valid(PENetwork_30_io_to_pes_21_in_valid),
    .io_to_pes_21_in_bits(PENetwork_30_io_to_pes_21_in_bits),
    .io_to_mem_valid(PENetwork_30_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_30_io_to_mem_bits)
  );
  PENetwork_22 PENetwork_31 ( // @[pe.scala 229:13]
    .io_to_pes_0_in_valid(PENetwork_31_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_31_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_31_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_31_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_31_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_31_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_31_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_31_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_31_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_31_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_31_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_31_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_31_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_31_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_31_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_31_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_31_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_31_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_31_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_31_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_31_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_31_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_31_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_31_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_31_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_31_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_31_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_31_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_31_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_31_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_31_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_31_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_31_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_31_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_31_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_31_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_31_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_31_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_31_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_31_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_31_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_31_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_31_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_31_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_31_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_31_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_31_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_31_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_31_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_31_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_31_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_31_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_31_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_31_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_31_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_31_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_31_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_31_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_31_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_31_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_31_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_31_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_31_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_31_io_to_pes_15_out_bits),
    .io_to_pes_16_in_valid(PENetwork_31_io_to_pes_16_in_valid),
    .io_to_pes_16_in_bits(PENetwork_31_io_to_pes_16_in_bits),
    .io_to_pes_16_out_valid(PENetwork_31_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_31_io_to_pes_16_out_bits),
    .io_to_pes_17_in_valid(PENetwork_31_io_to_pes_17_in_valid),
    .io_to_pes_17_in_bits(PENetwork_31_io_to_pes_17_in_bits),
    .io_to_pes_17_out_valid(PENetwork_31_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_31_io_to_pes_17_out_bits),
    .io_to_pes_18_in_valid(PENetwork_31_io_to_pes_18_in_valid),
    .io_to_pes_18_in_bits(PENetwork_31_io_to_pes_18_in_bits),
    .io_to_pes_18_out_valid(PENetwork_31_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_31_io_to_pes_18_out_bits),
    .io_to_pes_19_in_valid(PENetwork_31_io_to_pes_19_in_valid),
    .io_to_pes_19_in_bits(PENetwork_31_io_to_pes_19_in_bits),
    .io_to_pes_19_out_valid(PENetwork_31_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_31_io_to_pes_19_out_bits),
    .io_to_pes_20_in_valid(PENetwork_31_io_to_pes_20_in_valid),
    .io_to_pes_20_in_bits(PENetwork_31_io_to_pes_20_in_bits),
    .io_to_pes_20_out_valid(PENetwork_31_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_31_io_to_pes_20_out_bits),
    .io_to_pes_21_in_valid(PENetwork_31_io_to_pes_21_in_valid),
    .io_to_pes_21_in_bits(PENetwork_31_io_to_pes_21_in_bits),
    .io_to_mem_valid(PENetwork_31_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_31_io_to_mem_bits)
  );
  PENetwork_22 PENetwork_32 ( // @[pe.scala 229:13]
    .io_to_pes_0_in_valid(PENetwork_32_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_32_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_32_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_32_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_32_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_32_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_32_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_32_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_32_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_32_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_32_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_32_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_32_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_32_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_32_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_32_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_32_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_32_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_32_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_32_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_32_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_32_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_32_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_32_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_32_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_32_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_32_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_32_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_32_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_32_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_32_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_32_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_32_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_32_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_32_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_32_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_32_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_32_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_32_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_32_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_32_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_32_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_32_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_32_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_32_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_32_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_32_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_32_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_32_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_32_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_32_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_32_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_32_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_32_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_32_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_32_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_32_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_32_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_32_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_32_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_32_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_32_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_32_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_32_io_to_pes_15_out_bits),
    .io_to_pes_16_in_valid(PENetwork_32_io_to_pes_16_in_valid),
    .io_to_pes_16_in_bits(PENetwork_32_io_to_pes_16_in_bits),
    .io_to_pes_16_out_valid(PENetwork_32_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_32_io_to_pes_16_out_bits),
    .io_to_pes_17_in_valid(PENetwork_32_io_to_pes_17_in_valid),
    .io_to_pes_17_in_bits(PENetwork_32_io_to_pes_17_in_bits),
    .io_to_pes_17_out_valid(PENetwork_32_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_32_io_to_pes_17_out_bits),
    .io_to_pes_18_in_valid(PENetwork_32_io_to_pes_18_in_valid),
    .io_to_pes_18_in_bits(PENetwork_32_io_to_pes_18_in_bits),
    .io_to_pes_18_out_valid(PENetwork_32_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_32_io_to_pes_18_out_bits),
    .io_to_pes_19_in_valid(PENetwork_32_io_to_pes_19_in_valid),
    .io_to_pes_19_in_bits(PENetwork_32_io_to_pes_19_in_bits),
    .io_to_pes_19_out_valid(PENetwork_32_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_32_io_to_pes_19_out_bits),
    .io_to_pes_20_in_valid(PENetwork_32_io_to_pes_20_in_valid),
    .io_to_pes_20_in_bits(PENetwork_32_io_to_pes_20_in_bits),
    .io_to_pes_20_out_valid(PENetwork_32_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_32_io_to_pes_20_out_bits),
    .io_to_pes_21_in_valid(PENetwork_32_io_to_pes_21_in_valid),
    .io_to_pes_21_in_bits(PENetwork_32_io_to_pes_21_in_bits),
    .io_to_mem_valid(PENetwork_32_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_32_io_to_mem_bits)
  );
  PENetwork_22 PENetwork_33 ( // @[pe.scala 229:13]
    .io_to_pes_0_in_valid(PENetwork_33_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_33_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_33_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_33_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_33_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_33_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_33_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_33_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_33_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_33_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_33_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_33_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_33_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_33_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_33_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_33_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_33_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_33_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_33_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_33_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_33_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_33_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_33_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_33_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_33_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_33_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_33_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_33_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_33_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_33_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_33_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_33_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_33_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_33_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_33_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_33_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_33_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_33_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_33_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_33_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_33_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_33_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_33_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_33_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_33_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_33_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_33_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_33_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_33_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_33_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_33_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_33_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_33_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_33_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_33_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_33_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_33_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_33_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_33_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_33_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_33_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_33_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_33_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_33_io_to_pes_15_out_bits),
    .io_to_pes_16_in_valid(PENetwork_33_io_to_pes_16_in_valid),
    .io_to_pes_16_in_bits(PENetwork_33_io_to_pes_16_in_bits),
    .io_to_pes_16_out_valid(PENetwork_33_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_33_io_to_pes_16_out_bits),
    .io_to_pes_17_in_valid(PENetwork_33_io_to_pes_17_in_valid),
    .io_to_pes_17_in_bits(PENetwork_33_io_to_pes_17_in_bits),
    .io_to_pes_17_out_valid(PENetwork_33_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_33_io_to_pes_17_out_bits),
    .io_to_pes_18_in_valid(PENetwork_33_io_to_pes_18_in_valid),
    .io_to_pes_18_in_bits(PENetwork_33_io_to_pes_18_in_bits),
    .io_to_pes_18_out_valid(PENetwork_33_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_33_io_to_pes_18_out_bits),
    .io_to_pes_19_in_valid(PENetwork_33_io_to_pes_19_in_valid),
    .io_to_pes_19_in_bits(PENetwork_33_io_to_pes_19_in_bits),
    .io_to_pes_19_out_valid(PENetwork_33_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_33_io_to_pes_19_out_bits),
    .io_to_pes_20_in_valid(PENetwork_33_io_to_pes_20_in_valid),
    .io_to_pes_20_in_bits(PENetwork_33_io_to_pes_20_in_bits),
    .io_to_pes_20_out_valid(PENetwork_33_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_33_io_to_pes_20_out_bits),
    .io_to_pes_21_in_valid(PENetwork_33_io_to_pes_21_in_valid),
    .io_to_pes_21_in_bits(PENetwork_33_io_to_pes_21_in_bits),
    .io_to_mem_valid(PENetwork_33_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_33_io_to_mem_bits)
  );
  PENetwork_22 PENetwork_34 ( // @[pe.scala 229:13]
    .io_to_pes_0_in_valid(PENetwork_34_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_34_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_34_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_34_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_34_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_34_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_34_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_34_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_34_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_34_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_34_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_34_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_34_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_34_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_34_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_34_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_34_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_34_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_34_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_34_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_34_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_34_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_34_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_34_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_34_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_34_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_34_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_34_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_34_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_34_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_34_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_34_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_34_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_34_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_34_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_34_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_34_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_34_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_34_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_34_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_34_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_34_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_34_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_34_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_34_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_34_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_34_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_34_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_34_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_34_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_34_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_34_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_34_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_34_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_34_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_34_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_34_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_34_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_34_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_34_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_34_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_34_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_34_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_34_io_to_pes_15_out_bits),
    .io_to_pes_16_in_valid(PENetwork_34_io_to_pes_16_in_valid),
    .io_to_pes_16_in_bits(PENetwork_34_io_to_pes_16_in_bits),
    .io_to_pes_16_out_valid(PENetwork_34_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_34_io_to_pes_16_out_bits),
    .io_to_pes_17_in_valid(PENetwork_34_io_to_pes_17_in_valid),
    .io_to_pes_17_in_bits(PENetwork_34_io_to_pes_17_in_bits),
    .io_to_pes_17_out_valid(PENetwork_34_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_34_io_to_pes_17_out_bits),
    .io_to_pes_18_in_valid(PENetwork_34_io_to_pes_18_in_valid),
    .io_to_pes_18_in_bits(PENetwork_34_io_to_pes_18_in_bits),
    .io_to_pes_18_out_valid(PENetwork_34_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_34_io_to_pes_18_out_bits),
    .io_to_pes_19_in_valid(PENetwork_34_io_to_pes_19_in_valid),
    .io_to_pes_19_in_bits(PENetwork_34_io_to_pes_19_in_bits),
    .io_to_pes_19_out_valid(PENetwork_34_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_34_io_to_pes_19_out_bits),
    .io_to_pes_20_in_valid(PENetwork_34_io_to_pes_20_in_valid),
    .io_to_pes_20_in_bits(PENetwork_34_io_to_pes_20_in_bits),
    .io_to_pes_20_out_valid(PENetwork_34_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_34_io_to_pes_20_out_bits),
    .io_to_pes_21_in_valid(PENetwork_34_io_to_pes_21_in_valid),
    .io_to_pes_21_in_bits(PENetwork_34_io_to_pes_21_in_bits),
    .io_to_mem_valid(PENetwork_34_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_34_io_to_mem_bits)
  );
  PENetwork_22 PENetwork_35 ( // @[pe.scala 229:13]
    .io_to_pes_0_in_valid(PENetwork_35_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_35_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_35_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_35_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_35_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_35_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_35_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_35_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_35_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_35_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_35_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_35_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_35_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_35_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_35_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_35_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_35_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_35_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_35_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_35_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_35_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_35_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_35_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_35_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_35_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_35_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_35_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_35_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_35_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_35_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_35_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_35_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_35_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_35_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_35_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_35_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_35_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_35_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_35_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_35_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_35_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_35_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_35_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_35_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_35_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_35_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_35_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_35_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_35_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_35_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_35_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_35_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_35_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_35_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_35_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_35_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_35_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_35_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_35_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_35_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_35_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_35_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_35_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_35_io_to_pes_15_out_bits),
    .io_to_pes_16_in_valid(PENetwork_35_io_to_pes_16_in_valid),
    .io_to_pes_16_in_bits(PENetwork_35_io_to_pes_16_in_bits),
    .io_to_pes_16_out_valid(PENetwork_35_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_35_io_to_pes_16_out_bits),
    .io_to_pes_17_in_valid(PENetwork_35_io_to_pes_17_in_valid),
    .io_to_pes_17_in_bits(PENetwork_35_io_to_pes_17_in_bits),
    .io_to_pes_17_out_valid(PENetwork_35_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_35_io_to_pes_17_out_bits),
    .io_to_pes_18_in_valid(PENetwork_35_io_to_pes_18_in_valid),
    .io_to_pes_18_in_bits(PENetwork_35_io_to_pes_18_in_bits),
    .io_to_pes_18_out_valid(PENetwork_35_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_35_io_to_pes_18_out_bits),
    .io_to_pes_19_in_valid(PENetwork_35_io_to_pes_19_in_valid),
    .io_to_pes_19_in_bits(PENetwork_35_io_to_pes_19_in_bits),
    .io_to_pes_19_out_valid(PENetwork_35_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_35_io_to_pes_19_out_bits),
    .io_to_pes_20_in_valid(PENetwork_35_io_to_pes_20_in_valid),
    .io_to_pes_20_in_bits(PENetwork_35_io_to_pes_20_in_bits),
    .io_to_pes_20_out_valid(PENetwork_35_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_35_io_to_pes_20_out_bits),
    .io_to_pes_21_in_valid(PENetwork_35_io_to_pes_21_in_valid),
    .io_to_pes_21_in_bits(PENetwork_35_io_to_pes_21_in_bits),
    .io_to_mem_valid(PENetwork_35_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_35_io_to_mem_bits)
  );
  PENetwork_22 PENetwork_36 ( // @[pe.scala 229:13]
    .io_to_pes_0_in_valid(PENetwork_36_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_36_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_36_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_36_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_36_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_36_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_36_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_36_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_36_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_36_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_36_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_36_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_36_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_36_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_36_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_36_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_36_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_36_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_36_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_36_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_36_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_36_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_36_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_36_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_36_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_36_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_36_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_36_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_36_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_36_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_36_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_36_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_36_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_36_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_36_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_36_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_36_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_36_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_36_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_36_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_36_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_36_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_36_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_36_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_36_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_36_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_36_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_36_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_36_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_36_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_36_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_36_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_36_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_36_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_36_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_36_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_36_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_36_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_36_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_36_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_36_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_36_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_36_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_36_io_to_pes_15_out_bits),
    .io_to_pes_16_in_valid(PENetwork_36_io_to_pes_16_in_valid),
    .io_to_pes_16_in_bits(PENetwork_36_io_to_pes_16_in_bits),
    .io_to_pes_16_out_valid(PENetwork_36_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_36_io_to_pes_16_out_bits),
    .io_to_pes_17_in_valid(PENetwork_36_io_to_pes_17_in_valid),
    .io_to_pes_17_in_bits(PENetwork_36_io_to_pes_17_in_bits),
    .io_to_pes_17_out_valid(PENetwork_36_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_36_io_to_pes_17_out_bits),
    .io_to_pes_18_in_valid(PENetwork_36_io_to_pes_18_in_valid),
    .io_to_pes_18_in_bits(PENetwork_36_io_to_pes_18_in_bits),
    .io_to_pes_18_out_valid(PENetwork_36_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_36_io_to_pes_18_out_bits),
    .io_to_pes_19_in_valid(PENetwork_36_io_to_pes_19_in_valid),
    .io_to_pes_19_in_bits(PENetwork_36_io_to_pes_19_in_bits),
    .io_to_pes_19_out_valid(PENetwork_36_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_36_io_to_pes_19_out_bits),
    .io_to_pes_20_in_valid(PENetwork_36_io_to_pes_20_in_valid),
    .io_to_pes_20_in_bits(PENetwork_36_io_to_pes_20_in_bits),
    .io_to_pes_20_out_valid(PENetwork_36_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_36_io_to_pes_20_out_bits),
    .io_to_pes_21_in_valid(PENetwork_36_io_to_pes_21_in_valid),
    .io_to_pes_21_in_bits(PENetwork_36_io_to_pes_21_in_bits),
    .io_to_mem_valid(PENetwork_36_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_36_io_to_mem_bits)
  );
  PENetwork_22 PENetwork_37 ( // @[pe.scala 229:13]
    .io_to_pes_0_in_valid(PENetwork_37_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_37_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_37_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_37_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_37_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_37_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_37_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_37_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_37_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_37_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_37_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_37_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_37_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_37_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_37_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_37_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_37_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_37_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_37_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_37_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_37_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_37_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_37_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_37_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_37_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_37_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_37_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_37_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_37_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_37_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_37_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_37_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_37_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_37_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_37_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_37_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_37_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_37_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_37_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_37_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_37_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_37_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_37_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_37_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_37_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_37_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_37_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_37_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_37_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_37_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_37_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_37_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_37_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_37_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_37_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_37_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_37_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_37_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_37_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_37_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_37_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_37_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_37_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_37_io_to_pes_15_out_bits),
    .io_to_pes_16_in_valid(PENetwork_37_io_to_pes_16_in_valid),
    .io_to_pes_16_in_bits(PENetwork_37_io_to_pes_16_in_bits),
    .io_to_pes_16_out_valid(PENetwork_37_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_37_io_to_pes_16_out_bits),
    .io_to_pes_17_in_valid(PENetwork_37_io_to_pes_17_in_valid),
    .io_to_pes_17_in_bits(PENetwork_37_io_to_pes_17_in_bits),
    .io_to_pes_17_out_valid(PENetwork_37_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_37_io_to_pes_17_out_bits),
    .io_to_pes_18_in_valid(PENetwork_37_io_to_pes_18_in_valid),
    .io_to_pes_18_in_bits(PENetwork_37_io_to_pes_18_in_bits),
    .io_to_pes_18_out_valid(PENetwork_37_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_37_io_to_pes_18_out_bits),
    .io_to_pes_19_in_valid(PENetwork_37_io_to_pes_19_in_valid),
    .io_to_pes_19_in_bits(PENetwork_37_io_to_pes_19_in_bits),
    .io_to_pes_19_out_valid(PENetwork_37_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_37_io_to_pes_19_out_bits),
    .io_to_pes_20_in_valid(PENetwork_37_io_to_pes_20_in_valid),
    .io_to_pes_20_in_bits(PENetwork_37_io_to_pes_20_in_bits),
    .io_to_pes_20_out_valid(PENetwork_37_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_37_io_to_pes_20_out_bits),
    .io_to_pes_21_in_valid(PENetwork_37_io_to_pes_21_in_valid),
    .io_to_pes_21_in_bits(PENetwork_37_io_to_pes_21_in_bits),
    .io_to_mem_valid(PENetwork_37_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_37_io_to_mem_bits)
  );
  PENetwork_22 PENetwork_38 ( // @[pe.scala 229:13]
    .io_to_pes_0_in_valid(PENetwork_38_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_38_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_38_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_38_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_38_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_38_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_38_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_38_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_38_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_38_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_38_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_38_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_38_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_38_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_38_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_38_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_38_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_38_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_38_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_38_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_38_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_38_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_38_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_38_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_38_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_38_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_38_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_38_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_38_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_38_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_38_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_38_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_38_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_38_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_38_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_38_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_38_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_38_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_38_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_38_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_38_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_38_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_38_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_38_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_38_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_38_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_38_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_38_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_38_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_38_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_38_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_38_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_38_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_38_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_38_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_38_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_38_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_38_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_38_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_38_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_38_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_38_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_38_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_38_io_to_pes_15_out_bits),
    .io_to_pes_16_in_valid(PENetwork_38_io_to_pes_16_in_valid),
    .io_to_pes_16_in_bits(PENetwork_38_io_to_pes_16_in_bits),
    .io_to_pes_16_out_valid(PENetwork_38_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_38_io_to_pes_16_out_bits),
    .io_to_pes_17_in_valid(PENetwork_38_io_to_pes_17_in_valid),
    .io_to_pes_17_in_bits(PENetwork_38_io_to_pes_17_in_bits),
    .io_to_pes_17_out_valid(PENetwork_38_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_38_io_to_pes_17_out_bits),
    .io_to_pes_18_in_valid(PENetwork_38_io_to_pes_18_in_valid),
    .io_to_pes_18_in_bits(PENetwork_38_io_to_pes_18_in_bits),
    .io_to_pes_18_out_valid(PENetwork_38_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_38_io_to_pes_18_out_bits),
    .io_to_pes_19_in_valid(PENetwork_38_io_to_pes_19_in_valid),
    .io_to_pes_19_in_bits(PENetwork_38_io_to_pes_19_in_bits),
    .io_to_pes_19_out_valid(PENetwork_38_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_38_io_to_pes_19_out_bits),
    .io_to_pes_20_in_valid(PENetwork_38_io_to_pes_20_in_valid),
    .io_to_pes_20_in_bits(PENetwork_38_io_to_pes_20_in_bits),
    .io_to_pes_20_out_valid(PENetwork_38_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_38_io_to_pes_20_out_bits),
    .io_to_pes_21_in_valid(PENetwork_38_io_to_pes_21_in_valid),
    .io_to_pes_21_in_bits(PENetwork_38_io_to_pes_21_in_bits),
    .io_to_mem_valid(PENetwork_38_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_38_io_to_mem_bits)
  );
  PENetwork_22 PENetwork_39 ( // @[pe.scala 229:13]
    .io_to_pes_0_in_valid(PENetwork_39_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_39_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_39_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_39_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_39_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_39_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_39_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_39_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_39_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_39_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_39_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_39_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_39_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_39_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_39_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_39_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_39_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_39_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_39_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_39_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_39_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_39_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_39_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_39_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_39_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_39_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_39_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_39_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_39_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_39_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_39_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_39_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_39_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_39_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_39_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_39_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_39_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_39_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_39_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_39_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_39_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_39_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_39_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_39_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_39_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_39_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_39_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_39_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_39_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_39_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_39_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_39_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_39_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_39_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_39_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_39_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_39_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_39_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_39_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_39_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_39_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_39_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_39_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_39_io_to_pes_15_out_bits),
    .io_to_pes_16_in_valid(PENetwork_39_io_to_pes_16_in_valid),
    .io_to_pes_16_in_bits(PENetwork_39_io_to_pes_16_in_bits),
    .io_to_pes_16_out_valid(PENetwork_39_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_39_io_to_pes_16_out_bits),
    .io_to_pes_17_in_valid(PENetwork_39_io_to_pes_17_in_valid),
    .io_to_pes_17_in_bits(PENetwork_39_io_to_pes_17_in_bits),
    .io_to_pes_17_out_valid(PENetwork_39_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_39_io_to_pes_17_out_bits),
    .io_to_pes_18_in_valid(PENetwork_39_io_to_pes_18_in_valid),
    .io_to_pes_18_in_bits(PENetwork_39_io_to_pes_18_in_bits),
    .io_to_pes_18_out_valid(PENetwork_39_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_39_io_to_pes_18_out_bits),
    .io_to_pes_19_in_valid(PENetwork_39_io_to_pes_19_in_valid),
    .io_to_pes_19_in_bits(PENetwork_39_io_to_pes_19_in_bits),
    .io_to_pes_19_out_valid(PENetwork_39_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_39_io_to_pes_19_out_bits),
    .io_to_pes_20_in_valid(PENetwork_39_io_to_pes_20_in_valid),
    .io_to_pes_20_in_bits(PENetwork_39_io_to_pes_20_in_bits),
    .io_to_pes_20_out_valid(PENetwork_39_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_39_io_to_pes_20_out_bits),
    .io_to_pes_21_in_valid(PENetwork_39_io_to_pes_21_in_valid),
    .io_to_pes_21_in_bits(PENetwork_39_io_to_pes_21_in_bits),
    .io_to_mem_valid(PENetwork_39_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_39_io_to_mem_bits)
  );
  PENetwork_22 PENetwork_40 ( // @[pe.scala 229:13]
    .io_to_pes_0_in_valid(PENetwork_40_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_40_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_40_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_40_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_40_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_40_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_40_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_40_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_40_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_40_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_40_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_40_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_40_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_40_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_40_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_40_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_40_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_40_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_40_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_40_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_40_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_40_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_40_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_40_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_40_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_40_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_40_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_40_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_40_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_40_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_40_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_40_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_40_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_40_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_40_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_40_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_40_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_40_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_40_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_40_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_40_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_40_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_40_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_40_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_40_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_40_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_40_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_40_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_40_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_40_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_40_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_40_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_40_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_40_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_40_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_40_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_40_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_40_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_40_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_40_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_40_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_40_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_40_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_40_io_to_pes_15_out_bits),
    .io_to_pes_16_in_valid(PENetwork_40_io_to_pes_16_in_valid),
    .io_to_pes_16_in_bits(PENetwork_40_io_to_pes_16_in_bits),
    .io_to_pes_16_out_valid(PENetwork_40_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_40_io_to_pes_16_out_bits),
    .io_to_pes_17_in_valid(PENetwork_40_io_to_pes_17_in_valid),
    .io_to_pes_17_in_bits(PENetwork_40_io_to_pes_17_in_bits),
    .io_to_pes_17_out_valid(PENetwork_40_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_40_io_to_pes_17_out_bits),
    .io_to_pes_18_in_valid(PENetwork_40_io_to_pes_18_in_valid),
    .io_to_pes_18_in_bits(PENetwork_40_io_to_pes_18_in_bits),
    .io_to_pes_18_out_valid(PENetwork_40_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_40_io_to_pes_18_out_bits),
    .io_to_pes_19_in_valid(PENetwork_40_io_to_pes_19_in_valid),
    .io_to_pes_19_in_bits(PENetwork_40_io_to_pes_19_in_bits),
    .io_to_pes_19_out_valid(PENetwork_40_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_40_io_to_pes_19_out_bits),
    .io_to_pes_20_in_valid(PENetwork_40_io_to_pes_20_in_valid),
    .io_to_pes_20_in_bits(PENetwork_40_io_to_pes_20_in_bits),
    .io_to_pes_20_out_valid(PENetwork_40_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_40_io_to_pes_20_out_bits),
    .io_to_pes_21_in_valid(PENetwork_40_io_to_pes_21_in_valid),
    .io_to_pes_21_in_bits(PENetwork_40_io_to_pes_21_in_bits),
    .io_to_mem_valid(PENetwork_40_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_40_io_to_mem_bits)
  );
  PENetwork_22 PENetwork_41 ( // @[pe.scala 229:13]
    .io_to_pes_0_in_valid(PENetwork_41_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_41_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_41_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_41_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_41_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_41_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_41_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_41_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_41_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_41_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_41_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_41_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_41_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_41_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_41_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_41_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_41_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_41_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_41_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_41_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_41_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_41_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_41_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_41_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_41_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_41_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_41_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_41_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_41_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_41_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_41_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_41_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_41_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_41_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_41_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_41_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_41_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_41_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_41_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_41_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_41_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_41_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_41_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_41_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_41_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_41_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_41_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_41_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_41_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_41_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_41_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_41_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_41_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_41_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_41_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_41_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_41_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_41_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_41_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_41_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_41_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_41_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_41_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_41_io_to_pes_15_out_bits),
    .io_to_pes_16_in_valid(PENetwork_41_io_to_pes_16_in_valid),
    .io_to_pes_16_in_bits(PENetwork_41_io_to_pes_16_in_bits),
    .io_to_pes_16_out_valid(PENetwork_41_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_41_io_to_pes_16_out_bits),
    .io_to_pes_17_in_valid(PENetwork_41_io_to_pes_17_in_valid),
    .io_to_pes_17_in_bits(PENetwork_41_io_to_pes_17_in_bits),
    .io_to_pes_17_out_valid(PENetwork_41_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_41_io_to_pes_17_out_bits),
    .io_to_pes_18_in_valid(PENetwork_41_io_to_pes_18_in_valid),
    .io_to_pes_18_in_bits(PENetwork_41_io_to_pes_18_in_bits),
    .io_to_pes_18_out_valid(PENetwork_41_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_41_io_to_pes_18_out_bits),
    .io_to_pes_19_in_valid(PENetwork_41_io_to_pes_19_in_valid),
    .io_to_pes_19_in_bits(PENetwork_41_io_to_pes_19_in_bits),
    .io_to_pes_19_out_valid(PENetwork_41_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_41_io_to_pes_19_out_bits),
    .io_to_pes_20_in_valid(PENetwork_41_io_to_pes_20_in_valid),
    .io_to_pes_20_in_bits(PENetwork_41_io_to_pes_20_in_bits),
    .io_to_pes_20_out_valid(PENetwork_41_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_41_io_to_pes_20_out_bits),
    .io_to_pes_21_in_valid(PENetwork_41_io_to_pes_21_in_valid),
    .io_to_pes_21_in_bits(PENetwork_41_io_to_pes_21_in_bits),
    .io_to_mem_valid(PENetwork_41_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_41_io_to_mem_bits)
  );
  PENetwork_22 PENetwork_42 ( // @[pe.scala 229:13]
    .io_to_pes_0_in_valid(PENetwork_42_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_42_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_42_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_42_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_42_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_42_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_42_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_42_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_42_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_42_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_42_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_42_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_42_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_42_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_42_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_42_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_42_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_42_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_42_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_42_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_42_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_42_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_42_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_42_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_42_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_42_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_42_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_42_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_42_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_42_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_42_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_42_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_42_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_42_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_42_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_42_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_42_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_42_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_42_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_42_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_42_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_42_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_42_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_42_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_42_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_42_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_42_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_42_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_42_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_42_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_42_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_42_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_42_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_42_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_42_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_42_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_42_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_42_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_42_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_42_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_42_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_42_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_42_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_42_io_to_pes_15_out_bits),
    .io_to_pes_16_in_valid(PENetwork_42_io_to_pes_16_in_valid),
    .io_to_pes_16_in_bits(PENetwork_42_io_to_pes_16_in_bits),
    .io_to_pes_16_out_valid(PENetwork_42_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_42_io_to_pes_16_out_bits),
    .io_to_pes_17_in_valid(PENetwork_42_io_to_pes_17_in_valid),
    .io_to_pes_17_in_bits(PENetwork_42_io_to_pes_17_in_bits),
    .io_to_pes_17_out_valid(PENetwork_42_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_42_io_to_pes_17_out_bits),
    .io_to_pes_18_in_valid(PENetwork_42_io_to_pes_18_in_valid),
    .io_to_pes_18_in_bits(PENetwork_42_io_to_pes_18_in_bits),
    .io_to_pes_18_out_valid(PENetwork_42_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_42_io_to_pes_18_out_bits),
    .io_to_pes_19_in_valid(PENetwork_42_io_to_pes_19_in_valid),
    .io_to_pes_19_in_bits(PENetwork_42_io_to_pes_19_in_bits),
    .io_to_pes_19_out_valid(PENetwork_42_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_42_io_to_pes_19_out_bits),
    .io_to_pes_20_in_valid(PENetwork_42_io_to_pes_20_in_valid),
    .io_to_pes_20_in_bits(PENetwork_42_io_to_pes_20_in_bits),
    .io_to_pes_20_out_valid(PENetwork_42_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_42_io_to_pes_20_out_bits),
    .io_to_pes_21_in_valid(PENetwork_42_io_to_pes_21_in_valid),
    .io_to_pes_21_in_bits(PENetwork_42_io_to_pes_21_in_bits),
    .io_to_mem_valid(PENetwork_42_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_42_io_to_mem_bits)
  );
  PENetwork_22 PENetwork_43 ( // @[pe.scala 229:13]
    .io_to_pes_0_in_valid(PENetwork_43_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_43_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_43_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_43_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_43_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_43_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_43_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_43_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_43_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_43_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_43_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_43_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_43_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_43_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_43_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_43_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_43_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_43_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_43_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_43_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_43_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_43_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_43_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_43_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_43_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_43_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_43_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_43_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_43_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_43_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_43_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_43_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_43_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_43_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_43_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_43_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_43_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_43_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_43_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_43_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_43_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_43_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_43_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_43_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_43_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_43_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_43_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_43_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_43_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_43_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_43_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_43_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_43_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_43_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_43_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_43_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_43_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_43_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_43_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_43_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_43_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_43_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_43_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_43_io_to_pes_15_out_bits),
    .io_to_pes_16_in_valid(PENetwork_43_io_to_pes_16_in_valid),
    .io_to_pes_16_in_bits(PENetwork_43_io_to_pes_16_in_bits),
    .io_to_pes_16_out_valid(PENetwork_43_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_43_io_to_pes_16_out_bits),
    .io_to_pes_17_in_valid(PENetwork_43_io_to_pes_17_in_valid),
    .io_to_pes_17_in_bits(PENetwork_43_io_to_pes_17_in_bits),
    .io_to_pes_17_out_valid(PENetwork_43_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_43_io_to_pes_17_out_bits),
    .io_to_pes_18_in_valid(PENetwork_43_io_to_pes_18_in_valid),
    .io_to_pes_18_in_bits(PENetwork_43_io_to_pes_18_in_bits),
    .io_to_pes_18_out_valid(PENetwork_43_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_43_io_to_pes_18_out_bits),
    .io_to_pes_19_in_valid(PENetwork_43_io_to_pes_19_in_valid),
    .io_to_pes_19_in_bits(PENetwork_43_io_to_pes_19_in_bits),
    .io_to_pes_19_out_valid(PENetwork_43_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_43_io_to_pes_19_out_bits),
    .io_to_pes_20_in_valid(PENetwork_43_io_to_pes_20_in_valid),
    .io_to_pes_20_in_bits(PENetwork_43_io_to_pes_20_in_bits),
    .io_to_pes_20_out_valid(PENetwork_43_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_43_io_to_pes_20_out_bits),
    .io_to_pes_21_in_valid(PENetwork_43_io_to_pes_21_in_valid),
    .io_to_pes_21_in_bits(PENetwork_43_io_to_pes_21_in_bits),
    .io_to_mem_valid(PENetwork_43_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_43_io_to_mem_bits)
  );
  PENetwork_22 PENetwork_44 ( // @[pe.scala 229:13]
    .io_to_pes_0_in_valid(PENetwork_44_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_44_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_44_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_44_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_44_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_44_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_44_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_44_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_44_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_44_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_44_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_44_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_44_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_44_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_44_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_44_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_44_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_44_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_44_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_44_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_44_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_44_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_44_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_44_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_44_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_44_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_44_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_44_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_44_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_44_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_44_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_44_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_44_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_44_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_44_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_44_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_44_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_44_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_44_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_44_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_44_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_44_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_44_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_44_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_44_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_44_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_44_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_44_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_44_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_44_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_44_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_44_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_44_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_44_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_44_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_44_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_44_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_44_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_44_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_44_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_44_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_44_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_44_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_44_io_to_pes_15_out_bits),
    .io_to_pes_16_in_valid(PENetwork_44_io_to_pes_16_in_valid),
    .io_to_pes_16_in_bits(PENetwork_44_io_to_pes_16_in_bits),
    .io_to_pes_16_out_valid(PENetwork_44_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_44_io_to_pes_16_out_bits),
    .io_to_pes_17_in_valid(PENetwork_44_io_to_pes_17_in_valid),
    .io_to_pes_17_in_bits(PENetwork_44_io_to_pes_17_in_bits),
    .io_to_pes_17_out_valid(PENetwork_44_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_44_io_to_pes_17_out_bits),
    .io_to_pes_18_in_valid(PENetwork_44_io_to_pes_18_in_valid),
    .io_to_pes_18_in_bits(PENetwork_44_io_to_pes_18_in_bits),
    .io_to_pes_18_out_valid(PENetwork_44_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_44_io_to_pes_18_out_bits),
    .io_to_pes_19_in_valid(PENetwork_44_io_to_pes_19_in_valid),
    .io_to_pes_19_in_bits(PENetwork_44_io_to_pes_19_in_bits),
    .io_to_pes_19_out_valid(PENetwork_44_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_44_io_to_pes_19_out_bits),
    .io_to_pes_20_in_valid(PENetwork_44_io_to_pes_20_in_valid),
    .io_to_pes_20_in_bits(PENetwork_44_io_to_pes_20_in_bits),
    .io_to_pes_20_out_valid(PENetwork_44_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_44_io_to_pes_20_out_bits),
    .io_to_pes_21_in_valid(PENetwork_44_io_to_pes_21_in_valid),
    .io_to_pes_21_in_bits(PENetwork_44_io_to_pes_21_in_bits),
    .io_to_mem_valid(PENetwork_44_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_44_io_to_mem_bits)
  );
  PENetwork_22 PENetwork_45 ( // @[pe.scala 229:13]
    .io_to_pes_0_in_valid(PENetwork_45_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_45_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_45_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_45_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_45_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_45_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_45_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_45_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_45_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_45_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_45_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_45_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_45_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_45_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_45_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_45_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_45_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_45_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_45_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_45_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_45_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_45_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_45_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_45_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_45_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_45_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_45_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_45_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_45_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_45_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_45_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_45_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_45_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_45_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_45_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_45_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_45_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_45_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_45_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_45_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_45_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_45_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_45_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_45_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_45_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_45_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_45_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_45_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_45_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_45_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_45_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_45_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_45_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_45_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_45_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_45_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_45_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_45_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_45_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_45_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_45_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_45_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_45_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_45_io_to_pes_15_out_bits),
    .io_to_pes_16_in_valid(PENetwork_45_io_to_pes_16_in_valid),
    .io_to_pes_16_in_bits(PENetwork_45_io_to_pes_16_in_bits),
    .io_to_pes_16_out_valid(PENetwork_45_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_45_io_to_pes_16_out_bits),
    .io_to_pes_17_in_valid(PENetwork_45_io_to_pes_17_in_valid),
    .io_to_pes_17_in_bits(PENetwork_45_io_to_pes_17_in_bits),
    .io_to_pes_17_out_valid(PENetwork_45_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_45_io_to_pes_17_out_bits),
    .io_to_pes_18_in_valid(PENetwork_45_io_to_pes_18_in_valid),
    .io_to_pes_18_in_bits(PENetwork_45_io_to_pes_18_in_bits),
    .io_to_pes_18_out_valid(PENetwork_45_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_45_io_to_pes_18_out_bits),
    .io_to_pes_19_in_valid(PENetwork_45_io_to_pes_19_in_valid),
    .io_to_pes_19_in_bits(PENetwork_45_io_to_pes_19_in_bits),
    .io_to_pes_19_out_valid(PENetwork_45_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_45_io_to_pes_19_out_bits),
    .io_to_pes_20_in_valid(PENetwork_45_io_to_pes_20_in_valid),
    .io_to_pes_20_in_bits(PENetwork_45_io_to_pes_20_in_bits),
    .io_to_pes_20_out_valid(PENetwork_45_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_45_io_to_pes_20_out_bits),
    .io_to_pes_21_in_valid(PENetwork_45_io_to_pes_21_in_valid),
    .io_to_pes_21_in_bits(PENetwork_45_io_to_pes_21_in_bits),
    .io_to_mem_valid(PENetwork_45_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_45_io_to_mem_bits)
  );
  PENetwork_22 PENetwork_46 ( // @[pe.scala 229:13]
    .io_to_pes_0_in_valid(PENetwork_46_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_46_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_46_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_46_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_46_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_46_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_46_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_46_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_46_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_46_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_46_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_46_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_46_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_46_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_46_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_46_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_46_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_46_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_46_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_46_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_46_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_46_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_46_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_46_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_46_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_46_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_46_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_46_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_46_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_46_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_46_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_46_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_46_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_46_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_46_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_46_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_46_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_46_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_46_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_46_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_46_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_46_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_46_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_46_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_46_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_46_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_46_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_46_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_46_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_46_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_46_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_46_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_46_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_46_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_46_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_46_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_46_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_46_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_46_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_46_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_46_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_46_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_46_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_46_io_to_pes_15_out_bits),
    .io_to_pes_16_in_valid(PENetwork_46_io_to_pes_16_in_valid),
    .io_to_pes_16_in_bits(PENetwork_46_io_to_pes_16_in_bits),
    .io_to_pes_16_out_valid(PENetwork_46_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_46_io_to_pes_16_out_bits),
    .io_to_pes_17_in_valid(PENetwork_46_io_to_pes_17_in_valid),
    .io_to_pes_17_in_bits(PENetwork_46_io_to_pes_17_in_bits),
    .io_to_pes_17_out_valid(PENetwork_46_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_46_io_to_pes_17_out_bits),
    .io_to_pes_18_in_valid(PENetwork_46_io_to_pes_18_in_valid),
    .io_to_pes_18_in_bits(PENetwork_46_io_to_pes_18_in_bits),
    .io_to_pes_18_out_valid(PENetwork_46_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_46_io_to_pes_18_out_bits),
    .io_to_pes_19_in_valid(PENetwork_46_io_to_pes_19_in_valid),
    .io_to_pes_19_in_bits(PENetwork_46_io_to_pes_19_in_bits),
    .io_to_pes_19_out_valid(PENetwork_46_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_46_io_to_pes_19_out_bits),
    .io_to_pes_20_in_valid(PENetwork_46_io_to_pes_20_in_valid),
    .io_to_pes_20_in_bits(PENetwork_46_io_to_pes_20_in_bits),
    .io_to_pes_20_out_valid(PENetwork_46_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_46_io_to_pes_20_out_bits),
    .io_to_pes_21_in_valid(PENetwork_46_io_to_pes_21_in_valid),
    .io_to_pes_21_in_bits(PENetwork_46_io_to_pes_21_in_bits),
    .io_to_mem_valid(PENetwork_46_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_46_io_to_mem_bits)
  );
  PENetwork_22 PENetwork_47 ( // @[pe.scala 229:13]
    .io_to_pes_0_in_valid(PENetwork_47_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_47_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_47_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_47_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_47_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_47_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_47_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_47_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_47_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_47_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_47_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_47_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_47_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_47_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_47_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_47_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_47_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_47_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_47_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_47_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_47_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_47_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_47_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_47_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_47_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_47_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_47_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_47_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_47_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_47_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_47_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_47_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_47_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_47_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_47_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_47_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_47_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_47_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_47_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_47_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_47_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_47_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_47_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_47_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_47_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_47_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_47_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_47_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_47_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_47_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_47_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_47_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_47_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_47_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_47_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_47_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_47_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_47_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_47_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_47_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_47_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_47_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_47_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_47_io_to_pes_15_out_bits),
    .io_to_pes_16_in_valid(PENetwork_47_io_to_pes_16_in_valid),
    .io_to_pes_16_in_bits(PENetwork_47_io_to_pes_16_in_bits),
    .io_to_pes_16_out_valid(PENetwork_47_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_47_io_to_pes_16_out_bits),
    .io_to_pes_17_in_valid(PENetwork_47_io_to_pes_17_in_valid),
    .io_to_pes_17_in_bits(PENetwork_47_io_to_pes_17_in_bits),
    .io_to_pes_17_out_valid(PENetwork_47_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_47_io_to_pes_17_out_bits),
    .io_to_pes_18_in_valid(PENetwork_47_io_to_pes_18_in_valid),
    .io_to_pes_18_in_bits(PENetwork_47_io_to_pes_18_in_bits),
    .io_to_pes_18_out_valid(PENetwork_47_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_47_io_to_pes_18_out_bits),
    .io_to_pes_19_in_valid(PENetwork_47_io_to_pes_19_in_valid),
    .io_to_pes_19_in_bits(PENetwork_47_io_to_pes_19_in_bits),
    .io_to_pes_19_out_valid(PENetwork_47_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_47_io_to_pes_19_out_bits),
    .io_to_pes_20_in_valid(PENetwork_47_io_to_pes_20_in_valid),
    .io_to_pes_20_in_bits(PENetwork_47_io_to_pes_20_in_bits),
    .io_to_pes_20_out_valid(PENetwork_47_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_47_io_to_pes_20_out_bits),
    .io_to_pes_21_in_valid(PENetwork_47_io_to_pes_21_in_valid),
    .io_to_pes_21_in_bits(PENetwork_47_io_to_pes_21_in_bits),
    .io_to_mem_valid(PENetwork_47_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_47_io_to_mem_bits)
  );
  PENetwork_22 PENetwork_48 ( // @[pe.scala 229:13]
    .io_to_pes_0_in_valid(PENetwork_48_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_48_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_48_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_48_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_48_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_48_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_48_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_48_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_48_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_48_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_48_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_48_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_48_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_48_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_48_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_48_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_48_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_48_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_48_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_48_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_48_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_48_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_48_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_48_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_48_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_48_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_48_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_48_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_48_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_48_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_48_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_48_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_48_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_48_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_48_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_48_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_48_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_48_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_48_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_48_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_48_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_48_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_48_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_48_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_48_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_48_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_48_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_48_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_48_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_48_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_48_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_48_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_48_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_48_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_48_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_48_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_48_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_48_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_48_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_48_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_48_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_48_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_48_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_48_io_to_pes_15_out_bits),
    .io_to_pes_16_in_valid(PENetwork_48_io_to_pes_16_in_valid),
    .io_to_pes_16_in_bits(PENetwork_48_io_to_pes_16_in_bits),
    .io_to_pes_16_out_valid(PENetwork_48_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_48_io_to_pes_16_out_bits),
    .io_to_pes_17_in_valid(PENetwork_48_io_to_pes_17_in_valid),
    .io_to_pes_17_in_bits(PENetwork_48_io_to_pes_17_in_bits),
    .io_to_pes_17_out_valid(PENetwork_48_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_48_io_to_pes_17_out_bits),
    .io_to_pes_18_in_valid(PENetwork_48_io_to_pes_18_in_valid),
    .io_to_pes_18_in_bits(PENetwork_48_io_to_pes_18_in_bits),
    .io_to_pes_18_out_valid(PENetwork_48_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_48_io_to_pes_18_out_bits),
    .io_to_pes_19_in_valid(PENetwork_48_io_to_pes_19_in_valid),
    .io_to_pes_19_in_bits(PENetwork_48_io_to_pes_19_in_bits),
    .io_to_pes_19_out_valid(PENetwork_48_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_48_io_to_pes_19_out_bits),
    .io_to_pes_20_in_valid(PENetwork_48_io_to_pes_20_in_valid),
    .io_to_pes_20_in_bits(PENetwork_48_io_to_pes_20_in_bits),
    .io_to_pes_20_out_valid(PENetwork_48_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_48_io_to_pes_20_out_bits),
    .io_to_pes_21_in_valid(PENetwork_48_io_to_pes_21_in_valid),
    .io_to_pes_21_in_bits(PENetwork_48_io_to_pes_21_in_bits),
    .io_to_mem_valid(PENetwork_48_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_48_io_to_mem_bits)
  );
  PENetwork_22 PENetwork_49 ( // @[pe.scala 229:13]
    .io_to_pes_0_in_valid(PENetwork_49_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_49_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_49_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_49_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_49_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_49_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_49_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_49_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_49_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_49_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_49_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_49_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_49_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_49_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_49_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_49_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_49_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_49_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_49_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_49_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_49_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_49_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_49_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_49_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_49_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_49_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_49_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_49_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_49_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_49_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_49_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_49_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_49_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_49_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_49_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_49_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_49_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_49_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_49_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_49_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_49_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_49_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_49_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_49_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_49_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_49_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_49_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_49_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_49_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_49_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_49_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_49_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_49_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_49_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_49_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_49_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_49_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_49_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_49_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_49_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_49_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_49_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_49_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_49_io_to_pes_15_out_bits),
    .io_to_pes_16_in_valid(PENetwork_49_io_to_pes_16_in_valid),
    .io_to_pes_16_in_bits(PENetwork_49_io_to_pes_16_in_bits),
    .io_to_pes_16_out_valid(PENetwork_49_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_49_io_to_pes_16_out_bits),
    .io_to_pes_17_in_valid(PENetwork_49_io_to_pes_17_in_valid),
    .io_to_pes_17_in_bits(PENetwork_49_io_to_pes_17_in_bits),
    .io_to_pes_17_out_valid(PENetwork_49_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_49_io_to_pes_17_out_bits),
    .io_to_pes_18_in_valid(PENetwork_49_io_to_pes_18_in_valid),
    .io_to_pes_18_in_bits(PENetwork_49_io_to_pes_18_in_bits),
    .io_to_pes_18_out_valid(PENetwork_49_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_49_io_to_pes_18_out_bits),
    .io_to_pes_19_in_valid(PENetwork_49_io_to_pes_19_in_valid),
    .io_to_pes_19_in_bits(PENetwork_49_io_to_pes_19_in_bits),
    .io_to_pes_19_out_valid(PENetwork_49_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_49_io_to_pes_19_out_bits),
    .io_to_pes_20_in_valid(PENetwork_49_io_to_pes_20_in_valid),
    .io_to_pes_20_in_bits(PENetwork_49_io_to_pes_20_in_bits),
    .io_to_pes_20_out_valid(PENetwork_49_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_49_io_to_pes_20_out_bits),
    .io_to_pes_21_in_valid(PENetwork_49_io_to_pes_21_in_valid),
    .io_to_pes_21_in_bits(PENetwork_49_io_to_pes_21_in_bits),
    .io_to_mem_valid(PENetwork_49_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_49_io_to_mem_bits)
  );
  PENetwork_22 PENetwork_50 ( // @[pe.scala 229:13]
    .io_to_pes_0_in_valid(PENetwork_50_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_50_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_50_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_50_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_50_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_50_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_50_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_50_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_50_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_50_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_50_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_50_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_50_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_50_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_50_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_50_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_50_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_50_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_50_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_50_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_50_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_50_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_50_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_50_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_50_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_50_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_50_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_50_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_50_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_50_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_50_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_50_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_50_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_50_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_50_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_50_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_50_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_50_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_50_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_50_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_50_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_50_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_50_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_50_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_50_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_50_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_50_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_50_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_50_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_50_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_50_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_50_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_50_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_50_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_50_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_50_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_50_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_50_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_50_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_50_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_50_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_50_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_50_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_50_io_to_pes_15_out_bits),
    .io_to_pes_16_in_valid(PENetwork_50_io_to_pes_16_in_valid),
    .io_to_pes_16_in_bits(PENetwork_50_io_to_pes_16_in_bits),
    .io_to_pes_16_out_valid(PENetwork_50_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_50_io_to_pes_16_out_bits),
    .io_to_pes_17_in_valid(PENetwork_50_io_to_pes_17_in_valid),
    .io_to_pes_17_in_bits(PENetwork_50_io_to_pes_17_in_bits),
    .io_to_pes_17_out_valid(PENetwork_50_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_50_io_to_pes_17_out_bits),
    .io_to_pes_18_in_valid(PENetwork_50_io_to_pes_18_in_valid),
    .io_to_pes_18_in_bits(PENetwork_50_io_to_pes_18_in_bits),
    .io_to_pes_18_out_valid(PENetwork_50_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_50_io_to_pes_18_out_bits),
    .io_to_pes_19_in_valid(PENetwork_50_io_to_pes_19_in_valid),
    .io_to_pes_19_in_bits(PENetwork_50_io_to_pes_19_in_bits),
    .io_to_pes_19_out_valid(PENetwork_50_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_50_io_to_pes_19_out_bits),
    .io_to_pes_20_in_valid(PENetwork_50_io_to_pes_20_in_valid),
    .io_to_pes_20_in_bits(PENetwork_50_io_to_pes_20_in_bits),
    .io_to_pes_20_out_valid(PENetwork_50_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_50_io_to_pes_20_out_bits),
    .io_to_pes_21_in_valid(PENetwork_50_io_to_pes_21_in_valid),
    .io_to_pes_21_in_bits(PENetwork_50_io_to_pes_21_in_bits),
    .io_to_mem_valid(PENetwork_50_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_50_io_to_mem_bits)
  );
  PENetwork_22 PENetwork_51 ( // @[pe.scala 229:13]
    .io_to_pes_0_in_valid(PENetwork_51_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_51_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_51_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_51_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_51_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_51_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_51_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_51_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_51_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_51_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_51_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_51_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_51_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_51_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_51_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_51_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_51_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_51_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_51_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_51_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_51_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_51_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_51_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_51_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_51_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_51_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_51_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_51_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_51_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_51_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_51_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_51_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_51_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_51_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_51_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_51_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_51_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_51_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_51_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_51_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_51_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_51_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_51_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_51_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_51_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_51_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_51_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_51_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_51_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_51_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_51_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_51_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_51_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_51_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_51_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_51_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_51_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_51_io_to_pes_14_in_bits),
    .io_to_pes_14_out_valid(PENetwork_51_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_51_io_to_pes_14_out_bits),
    .io_to_pes_15_in_valid(PENetwork_51_io_to_pes_15_in_valid),
    .io_to_pes_15_in_bits(PENetwork_51_io_to_pes_15_in_bits),
    .io_to_pes_15_out_valid(PENetwork_51_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_51_io_to_pes_15_out_bits),
    .io_to_pes_16_in_valid(PENetwork_51_io_to_pes_16_in_valid),
    .io_to_pes_16_in_bits(PENetwork_51_io_to_pes_16_in_bits),
    .io_to_pes_16_out_valid(PENetwork_51_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_51_io_to_pes_16_out_bits),
    .io_to_pes_17_in_valid(PENetwork_51_io_to_pes_17_in_valid),
    .io_to_pes_17_in_bits(PENetwork_51_io_to_pes_17_in_bits),
    .io_to_pes_17_out_valid(PENetwork_51_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_51_io_to_pes_17_out_bits),
    .io_to_pes_18_in_valid(PENetwork_51_io_to_pes_18_in_valid),
    .io_to_pes_18_in_bits(PENetwork_51_io_to_pes_18_in_bits),
    .io_to_pes_18_out_valid(PENetwork_51_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_51_io_to_pes_18_out_bits),
    .io_to_pes_19_in_valid(PENetwork_51_io_to_pes_19_in_valid),
    .io_to_pes_19_in_bits(PENetwork_51_io_to_pes_19_in_bits),
    .io_to_pes_19_out_valid(PENetwork_51_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_51_io_to_pes_19_out_bits),
    .io_to_pes_20_in_valid(PENetwork_51_io_to_pes_20_in_valid),
    .io_to_pes_20_in_bits(PENetwork_51_io_to_pes_20_in_bits),
    .io_to_pes_20_out_valid(PENetwork_51_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_51_io_to_pes_20_out_bits),
    .io_to_pes_21_in_valid(PENetwork_51_io_to_pes_21_in_valid),
    .io_to_pes_21_in_bits(PENetwork_51_io_to_pes_21_in_bits),
    .io_to_mem_valid(PENetwork_51_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_51_io_to_mem_bits)
  );
  PENetwork_52 PENetwork_52 ( // @[pe.scala 229:13]
    .clock(PENetwork_52_clock),
    .reset(PENetwork_52_reset),
    .io_to_pes_0_out_valid(PENetwork_52_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_52_io_to_pes_0_out_bits),
    .io_to_pes_0_sig_stat2trans(PENetwork_52_io_to_pes_0_sig_stat2trans),
    .io_to_pes_1_out_valid(PENetwork_52_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_52_io_to_pes_1_out_bits),
    .io_to_pes_1_sig_stat2trans(PENetwork_52_io_to_pes_1_sig_stat2trans),
    .io_to_pes_2_out_valid(PENetwork_52_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_52_io_to_pes_2_out_bits),
    .io_to_pes_2_sig_stat2trans(PENetwork_52_io_to_pes_2_sig_stat2trans),
    .io_to_pes_3_out_valid(PENetwork_52_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_52_io_to_pes_3_out_bits),
    .io_to_pes_3_sig_stat2trans(PENetwork_52_io_to_pes_3_sig_stat2trans),
    .io_to_pes_4_out_valid(PENetwork_52_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_52_io_to_pes_4_out_bits),
    .io_to_pes_4_sig_stat2trans(PENetwork_52_io_to_pes_4_sig_stat2trans),
    .io_to_pes_5_out_valid(PENetwork_52_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_52_io_to_pes_5_out_bits),
    .io_to_pes_5_sig_stat2trans(PENetwork_52_io_to_pes_5_sig_stat2trans),
    .io_to_pes_6_out_valid(PENetwork_52_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_52_io_to_pes_6_out_bits),
    .io_to_pes_6_sig_stat2trans(PENetwork_52_io_to_pes_6_sig_stat2trans),
    .io_to_pes_7_out_valid(PENetwork_52_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_52_io_to_pes_7_out_bits),
    .io_to_pes_7_sig_stat2trans(PENetwork_52_io_to_pes_7_sig_stat2trans),
    .io_to_pes_8_out_valid(PENetwork_52_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_52_io_to_pes_8_out_bits),
    .io_to_pes_8_sig_stat2trans(PENetwork_52_io_to_pes_8_sig_stat2trans),
    .io_to_pes_9_out_valid(PENetwork_52_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_52_io_to_pes_9_out_bits),
    .io_to_pes_9_sig_stat2trans(PENetwork_52_io_to_pes_9_sig_stat2trans),
    .io_to_pes_10_out_valid(PENetwork_52_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_52_io_to_pes_10_out_bits),
    .io_to_pes_10_sig_stat2trans(PENetwork_52_io_to_pes_10_sig_stat2trans),
    .io_to_pes_11_out_valid(PENetwork_52_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_52_io_to_pes_11_out_bits),
    .io_to_pes_11_sig_stat2trans(PENetwork_52_io_to_pes_11_sig_stat2trans),
    .io_to_pes_12_out_valid(PENetwork_52_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_52_io_to_pes_12_out_bits),
    .io_to_pes_12_sig_stat2trans(PENetwork_52_io_to_pes_12_sig_stat2trans),
    .io_to_pes_13_out_valid(PENetwork_52_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_52_io_to_pes_13_out_bits),
    .io_to_pes_13_sig_stat2trans(PENetwork_52_io_to_pes_13_sig_stat2trans),
    .io_to_pes_14_out_valid(PENetwork_52_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_52_io_to_pes_14_out_bits),
    .io_to_pes_14_sig_stat2trans(PENetwork_52_io_to_pes_14_sig_stat2trans),
    .io_to_pes_15_out_valid(PENetwork_52_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_52_io_to_pes_15_out_bits),
    .io_to_pes_15_sig_stat2trans(PENetwork_52_io_to_pes_15_sig_stat2trans),
    .io_to_pes_16_out_valid(PENetwork_52_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_52_io_to_pes_16_out_bits),
    .io_to_pes_16_sig_stat2trans(PENetwork_52_io_to_pes_16_sig_stat2trans),
    .io_to_pes_17_out_valid(PENetwork_52_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_52_io_to_pes_17_out_bits),
    .io_to_pes_17_sig_stat2trans(PENetwork_52_io_to_pes_17_sig_stat2trans),
    .io_to_pes_18_out_valid(PENetwork_52_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_52_io_to_pes_18_out_bits),
    .io_to_pes_18_sig_stat2trans(PENetwork_52_io_to_pes_18_sig_stat2trans),
    .io_to_pes_19_out_valid(PENetwork_52_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_52_io_to_pes_19_out_bits),
    .io_to_pes_19_sig_stat2trans(PENetwork_52_io_to_pes_19_sig_stat2trans),
    .io_to_pes_20_out_valid(PENetwork_52_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_52_io_to_pes_20_out_bits),
    .io_to_pes_20_sig_stat2trans(PENetwork_52_io_to_pes_20_sig_stat2trans),
    .io_to_pes_21_out_valid(PENetwork_52_io_to_pes_21_out_valid),
    .io_to_pes_21_out_bits(PENetwork_52_io_to_pes_21_out_bits),
    .io_to_pes_21_sig_stat2trans(PENetwork_52_io_to_pes_21_sig_stat2trans),
    .io_to_mem_valid(PENetwork_52_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_52_io_to_mem_bits),
    .io_sig_stat2trans(PENetwork_52_io_sig_stat2trans)
  );
  PENetwork_52 PENetwork_53 ( // @[pe.scala 229:13]
    .clock(PENetwork_53_clock),
    .reset(PENetwork_53_reset),
    .io_to_pes_0_out_valid(PENetwork_53_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_53_io_to_pes_0_out_bits),
    .io_to_pes_0_sig_stat2trans(PENetwork_53_io_to_pes_0_sig_stat2trans),
    .io_to_pes_1_out_valid(PENetwork_53_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_53_io_to_pes_1_out_bits),
    .io_to_pes_1_sig_stat2trans(PENetwork_53_io_to_pes_1_sig_stat2trans),
    .io_to_pes_2_out_valid(PENetwork_53_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_53_io_to_pes_2_out_bits),
    .io_to_pes_2_sig_stat2trans(PENetwork_53_io_to_pes_2_sig_stat2trans),
    .io_to_pes_3_out_valid(PENetwork_53_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_53_io_to_pes_3_out_bits),
    .io_to_pes_3_sig_stat2trans(PENetwork_53_io_to_pes_3_sig_stat2trans),
    .io_to_pes_4_out_valid(PENetwork_53_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_53_io_to_pes_4_out_bits),
    .io_to_pes_4_sig_stat2trans(PENetwork_53_io_to_pes_4_sig_stat2trans),
    .io_to_pes_5_out_valid(PENetwork_53_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_53_io_to_pes_5_out_bits),
    .io_to_pes_5_sig_stat2trans(PENetwork_53_io_to_pes_5_sig_stat2trans),
    .io_to_pes_6_out_valid(PENetwork_53_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_53_io_to_pes_6_out_bits),
    .io_to_pes_6_sig_stat2trans(PENetwork_53_io_to_pes_6_sig_stat2trans),
    .io_to_pes_7_out_valid(PENetwork_53_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_53_io_to_pes_7_out_bits),
    .io_to_pes_7_sig_stat2trans(PENetwork_53_io_to_pes_7_sig_stat2trans),
    .io_to_pes_8_out_valid(PENetwork_53_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_53_io_to_pes_8_out_bits),
    .io_to_pes_8_sig_stat2trans(PENetwork_53_io_to_pes_8_sig_stat2trans),
    .io_to_pes_9_out_valid(PENetwork_53_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_53_io_to_pes_9_out_bits),
    .io_to_pes_9_sig_stat2trans(PENetwork_53_io_to_pes_9_sig_stat2trans),
    .io_to_pes_10_out_valid(PENetwork_53_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_53_io_to_pes_10_out_bits),
    .io_to_pes_10_sig_stat2trans(PENetwork_53_io_to_pes_10_sig_stat2trans),
    .io_to_pes_11_out_valid(PENetwork_53_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_53_io_to_pes_11_out_bits),
    .io_to_pes_11_sig_stat2trans(PENetwork_53_io_to_pes_11_sig_stat2trans),
    .io_to_pes_12_out_valid(PENetwork_53_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_53_io_to_pes_12_out_bits),
    .io_to_pes_12_sig_stat2trans(PENetwork_53_io_to_pes_12_sig_stat2trans),
    .io_to_pes_13_out_valid(PENetwork_53_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_53_io_to_pes_13_out_bits),
    .io_to_pes_13_sig_stat2trans(PENetwork_53_io_to_pes_13_sig_stat2trans),
    .io_to_pes_14_out_valid(PENetwork_53_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_53_io_to_pes_14_out_bits),
    .io_to_pes_14_sig_stat2trans(PENetwork_53_io_to_pes_14_sig_stat2trans),
    .io_to_pes_15_out_valid(PENetwork_53_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_53_io_to_pes_15_out_bits),
    .io_to_pes_15_sig_stat2trans(PENetwork_53_io_to_pes_15_sig_stat2trans),
    .io_to_pes_16_out_valid(PENetwork_53_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_53_io_to_pes_16_out_bits),
    .io_to_pes_16_sig_stat2trans(PENetwork_53_io_to_pes_16_sig_stat2trans),
    .io_to_pes_17_out_valid(PENetwork_53_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_53_io_to_pes_17_out_bits),
    .io_to_pes_17_sig_stat2trans(PENetwork_53_io_to_pes_17_sig_stat2trans),
    .io_to_pes_18_out_valid(PENetwork_53_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_53_io_to_pes_18_out_bits),
    .io_to_pes_18_sig_stat2trans(PENetwork_53_io_to_pes_18_sig_stat2trans),
    .io_to_pes_19_out_valid(PENetwork_53_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_53_io_to_pes_19_out_bits),
    .io_to_pes_19_sig_stat2trans(PENetwork_53_io_to_pes_19_sig_stat2trans),
    .io_to_pes_20_out_valid(PENetwork_53_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_53_io_to_pes_20_out_bits),
    .io_to_pes_20_sig_stat2trans(PENetwork_53_io_to_pes_20_sig_stat2trans),
    .io_to_pes_21_out_valid(PENetwork_53_io_to_pes_21_out_valid),
    .io_to_pes_21_out_bits(PENetwork_53_io_to_pes_21_out_bits),
    .io_to_pes_21_sig_stat2trans(PENetwork_53_io_to_pes_21_sig_stat2trans),
    .io_to_mem_valid(PENetwork_53_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_53_io_to_mem_bits),
    .io_sig_stat2trans(PENetwork_53_io_sig_stat2trans)
  );
  PENetwork_52 PENetwork_54 ( // @[pe.scala 229:13]
    .clock(PENetwork_54_clock),
    .reset(PENetwork_54_reset),
    .io_to_pes_0_out_valid(PENetwork_54_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_54_io_to_pes_0_out_bits),
    .io_to_pes_0_sig_stat2trans(PENetwork_54_io_to_pes_0_sig_stat2trans),
    .io_to_pes_1_out_valid(PENetwork_54_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_54_io_to_pes_1_out_bits),
    .io_to_pes_1_sig_stat2trans(PENetwork_54_io_to_pes_1_sig_stat2trans),
    .io_to_pes_2_out_valid(PENetwork_54_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_54_io_to_pes_2_out_bits),
    .io_to_pes_2_sig_stat2trans(PENetwork_54_io_to_pes_2_sig_stat2trans),
    .io_to_pes_3_out_valid(PENetwork_54_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_54_io_to_pes_3_out_bits),
    .io_to_pes_3_sig_stat2trans(PENetwork_54_io_to_pes_3_sig_stat2trans),
    .io_to_pes_4_out_valid(PENetwork_54_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_54_io_to_pes_4_out_bits),
    .io_to_pes_4_sig_stat2trans(PENetwork_54_io_to_pes_4_sig_stat2trans),
    .io_to_pes_5_out_valid(PENetwork_54_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_54_io_to_pes_5_out_bits),
    .io_to_pes_5_sig_stat2trans(PENetwork_54_io_to_pes_5_sig_stat2trans),
    .io_to_pes_6_out_valid(PENetwork_54_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_54_io_to_pes_6_out_bits),
    .io_to_pes_6_sig_stat2trans(PENetwork_54_io_to_pes_6_sig_stat2trans),
    .io_to_pes_7_out_valid(PENetwork_54_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_54_io_to_pes_7_out_bits),
    .io_to_pes_7_sig_stat2trans(PENetwork_54_io_to_pes_7_sig_stat2trans),
    .io_to_pes_8_out_valid(PENetwork_54_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_54_io_to_pes_8_out_bits),
    .io_to_pes_8_sig_stat2trans(PENetwork_54_io_to_pes_8_sig_stat2trans),
    .io_to_pes_9_out_valid(PENetwork_54_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_54_io_to_pes_9_out_bits),
    .io_to_pes_9_sig_stat2trans(PENetwork_54_io_to_pes_9_sig_stat2trans),
    .io_to_pes_10_out_valid(PENetwork_54_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_54_io_to_pes_10_out_bits),
    .io_to_pes_10_sig_stat2trans(PENetwork_54_io_to_pes_10_sig_stat2trans),
    .io_to_pes_11_out_valid(PENetwork_54_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_54_io_to_pes_11_out_bits),
    .io_to_pes_11_sig_stat2trans(PENetwork_54_io_to_pes_11_sig_stat2trans),
    .io_to_pes_12_out_valid(PENetwork_54_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_54_io_to_pes_12_out_bits),
    .io_to_pes_12_sig_stat2trans(PENetwork_54_io_to_pes_12_sig_stat2trans),
    .io_to_pes_13_out_valid(PENetwork_54_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_54_io_to_pes_13_out_bits),
    .io_to_pes_13_sig_stat2trans(PENetwork_54_io_to_pes_13_sig_stat2trans),
    .io_to_pes_14_out_valid(PENetwork_54_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_54_io_to_pes_14_out_bits),
    .io_to_pes_14_sig_stat2trans(PENetwork_54_io_to_pes_14_sig_stat2trans),
    .io_to_pes_15_out_valid(PENetwork_54_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_54_io_to_pes_15_out_bits),
    .io_to_pes_15_sig_stat2trans(PENetwork_54_io_to_pes_15_sig_stat2trans),
    .io_to_pes_16_out_valid(PENetwork_54_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_54_io_to_pes_16_out_bits),
    .io_to_pes_16_sig_stat2trans(PENetwork_54_io_to_pes_16_sig_stat2trans),
    .io_to_pes_17_out_valid(PENetwork_54_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_54_io_to_pes_17_out_bits),
    .io_to_pes_17_sig_stat2trans(PENetwork_54_io_to_pes_17_sig_stat2trans),
    .io_to_pes_18_out_valid(PENetwork_54_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_54_io_to_pes_18_out_bits),
    .io_to_pes_18_sig_stat2trans(PENetwork_54_io_to_pes_18_sig_stat2trans),
    .io_to_pes_19_out_valid(PENetwork_54_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_54_io_to_pes_19_out_bits),
    .io_to_pes_19_sig_stat2trans(PENetwork_54_io_to_pes_19_sig_stat2trans),
    .io_to_pes_20_out_valid(PENetwork_54_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_54_io_to_pes_20_out_bits),
    .io_to_pes_20_sig_stat2trans(PENetwork_54_io_to_pes_20_sig_stat2trans),
    .io_to_pes_21_out_valid(PENetwork_54_io_to_pes_21_out_valid),
    .io_to_pes_21_out_bits(PENetwork_54_io_to_pes_21_out_bits),
    .io_to_pes_21_sig_stat2trans(PENetwork_54_io_to_pes_21_sig_stat2trans),
    .io_to_mem_valid(PENetwork_54_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_54_io_to_mem_bits),
    .io_sig_stat2trans(PENetwork_54_io_sig_stat2trans)
  );
  PENetwork_52 PENetwork_55 ( // @[pe.scala 229:13]
    .clock(PENetwork_55_clock),
    .reset(PENetwork_55_reset),
    .io_to_pes_0_out_valid(PENetwork_55_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_55_io_to_pes_0_out_bits),
    .io_to_pes_0_sig_stat2trans(PENetwork_55_io_to_pes_0_sig_stat2trans),
    .io_to_pes_1_out_valid(PENetwork_55_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_55_io_to_pes_1_out_bits),
    .io_to_pes_1_sig_stat2trans(PENetwork_55_io_to_pes_1_sig_stat2trans),
    .io_to_pes_2_out_valid(PENetwork_55_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_55_io_to_pes_2_out_bits),
    .io_to_pes_2_sig_stat2trans(PENetwork_55_io_to_pes_2_sig_stat2trans),
    .io_to_pes_3_out_valid(PENetwork_55_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_55_io_to_pes_3_out_bits),
    .io_to_pes_3_sig_stat2trans(PENetwork_55_io_to_pes_3_sig_stat2trans),
    .io_to_pes_4_out_valid(PENetwork_55_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_55_io_to_pes_4_out_bits),
    .io_to_pes_4_sig_stat2trans(PENetwork_55_io_to_pes_4_sig_stat2trans),
    .io_to_pes_5_out_valid(PENetwork_55_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_55_io_to_pes_5_out_bits),
    .io_to_pes_5_sig_stat2trans(PENetwork_55_io_to_pes_5_sig_stat2trans),
    .io_to_pes_6_out_valid(PENetwork_55_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_55_io_to_pes_6_out_bits),
    .io_to_pes_6_sig_stat2trans(PENetwork_55_io_to_pes_6_sig_stat2trans),
    .io_to_pes_7_out_valid(PENetwork_55_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_55_io_to_pes_7_out_bits),
    .io_to_pes_7_sig_stat2trans(PENetwork_55_io_to_pes_7_sig_stat2trans),
    .io_to_pes_8_out_valid(PENetwork_55_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_55_io_to_pes_8_out_bits),
    .io_to_pes_8_sig_stat2trans(PENetwork_55_io_to_pes_8_sig_stat2trans),
    .io_to_pes_9_out_valid(PENetwork_55_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_55_io_to_pes_9_out_bits),
    .io_to_pes_9_sig_stat2trans(PENetwork_55_io_to_pes_9_sig_stat2trans),
    .io_to_pes_10_out_valid(PENetwork_55_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_55_io_to_pes_10_out_bits),
    .io_to_pes_10_sig_stat2trans(PENetwork_55_io_to_pes_10_sig_stat2trans),
    .io_to_pes_11_out_valid(PENetwork_55_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_55_io_to_pes_11_out_bits),
    .io_to_pes_11_sig_stat2trans(PENetwork_55_io_to_pes_11_sig_stat2trans),
    .io_to_pes_12_out_valid(PENetwork_55_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_55_io_to_pes_12_out_bits),
    .io_to_pes_12_sig_stat2trans(PENetwork_55_io_to_pes_12_sig_stat2trans),
    .io_to_pes_13_out_valid(PENetwork_55_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_55_io_to_pes_13_out_bits),
    .io_to_pes_13_sig_stat2trans(PENetwork_55_io_to_pes_13_sig_stat2trans),
    .io_to_pes_14_out_valid(PENetwork_55_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_55_io_to_pes_14_out_bits),
    .io_to_pes_14_sig_stat2trans(PENetwork_55_io_to_pes_14_sig_stat2trans),
    .io_to_pes_15_out_valid(PENetwork_55_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_55_io_to_pes_15_out_bits),
    .io_to_pes_15_sig_stat2trans(PENetwork_55_io_to_pes_15_sig_stat2trans),
    .io_to_pes_16_out_valid(PENetwork_55_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_55_io_to_pes_16_out_bits),
    .io_to_pes_16_sig_stat2trans(PENetwork_55_io_to_pes_16_sig_stat2trans),
    .io_to_pes_17_out_valid(PENetwork_55_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_55_io_to_pes_17_out_bits),
    .io_to_pes_17_sig_stat2trans(PENetwork_55_io_to_pes_17_sig_stat2trans),
    .io_to_pes_18_out_valid(PENetwork_55_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_55_io_to_pes_18_out_bits),
    .io_to_pes_18_sig_stat2trans(PENetwork_55_io_to_pes_18_sig_stat2trans),
    .io_to_pes_19_out_valid(PENetwork_55_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_55_io_to_pes_19_out_bits),
    .io_to_pes_19_sig_stat2trans(PENetwork_55_io_to_pes_19_sig_stat2trans),
    .io_to_pes_20_out_valid(PENetwork_55_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_55_io_to_pes_20_out_bits),
    .io_to_pes_20_sig_stat2trans(PENetwork_55_io_to_pes_20_sig_stat2trans),
    .io_to_pes_21_out_valid(PENetwork_55_io_to_pes_21_out_valid),
    .io_to_pes_21_out_bits(PENetwork_55_io_to_pes_21_out_bits),
    .io_to_pes_21_sig_stat2trans(PENetwork_55_io_to_pes_21_sig_stat2trans),
    .io_to_mem_valid(PENetwork_55_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_55_io_to_mem_bits),
    .io_sig_stat2trans(PENetwork_55_io_sig_stat2trans)
  );
  PENetwork_52 PENetwork_56 ( // @[pe.scala 229:13]
    .clock(PENetwork_56_clock),
    .reset(PENetwork_56_reset),
    .io_to_pes_0_out_valid(PENetwork_56_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_56_io_to_pes_0_out_bits),
    .io_to_pes_0_sig_stat2trans(PENetwork_56_io_to_pes_0_sig_stat2trans),
    .io_to_pes_1_out_valid(PENetwork_56_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_56_io_to_pes_1_out_bits),
    .io_to_pes_1_sig_stat2trans(PENetwork_56_io_to_pes_1_sig_stat2trans),
    .io_to_pes_2_out_valid(PENetwork_56_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_56_io_to_pes_2_out_bits),
    .io_to_pes_2_sig_stat2trans(PENetwork_56_io_to_pes_2_sig_stat2trans),
    .io_to_pes_3_out_valid(PENetwork_56_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_56_io_to_pes_3_out_bits),
    .io_to_pes_3_sig_stat2trans(PENetwork_56_io_to_pes_3_sig_stat2trans),
    .io_to_pes_4_out_valid(PENetwork_56_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_56_io_to_pes_4_out_bits),
    .io_to_pes_4_sig_stat2trans(PENetwork_56_io_to_pes_4_sig_stat2trans),
    .io_to_pes_5_out_valid(PENetwork_56_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_56_io_to_pes_5_out_bits),
    .io_to_pes_5_sig_stat2trans(PENetwork_56_io_to_pes_5_sig_stat2trans),
    .io_to_pes_6_out_valid(PENetwork_56_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_56_io_to_pes_6_out_bits),
    .io_to_pes_6_sig_stat2trans(PENetwork_56_io_to_pes_6_sig_stat2trans),
    .io_to_pes_7_out_valid(PENetwork_56_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_56_io_to_pes_7_out_bits),
    .io_to_pes_7_sig_stat2trans(PENetwork_56_io_to_pes_7_sig_stat2trans),
    .io_to_pes_8_out_valid(PENetwork_56_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_56_io_to_pes_8_out_bits),
    .io_to_pes_8_sig_stat2trans(PENetwork_56_io_to_pes_8_sig_stat2trans),
    .io_to_pes_9_out_valid(PENetwork_56_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_56_io_to_pes_9_out_bits),
    .io_to_pes_9_sig_stat2trans(PENetwork_56_io_to_pes_9_sig_stat2trans),
    .io_to_pes_10_out_valid(PENetwork_56_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_56_io_to_pes_10_out_bits),
    .io_to_pes_10_sig_stat2trans(PENetwork_56_io_to_pes_10_sig_stat2trans),
    .io_to_pes_11_out_valid(PENetwork_56_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_56_io_to_pes_11_out_bits),
    .io_to_pes_11_sig_stat2trans(PENetwork_56_io_to_pes_11_sig_stat2trans),
    .io_to_pes_12_out_valid(PENetwork_56_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_56_io_to_pes_12_out_bits),
    .io_to_pes_12_sig_stat2trans(PENetwork_56_io_to_pes_12_sig_stat2trans),
    .io_to_pes_13_out_valid(PENetwork_56_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_56_io_to_pes_13_out_bits),
    .io_to_pes_13_sig_stat2trans(PENetwork_56_io_to_pes_13_sig_stat2trans),
    .io_to_pes_14_out_valid(PENetwork_56_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_56_io_to_pes_14_out_bits),
    .io_to_pes_14_sig_stat2trans(PENetwork_56_io_to_pes_14_sig_stat2trans),
    .io_to_pes_15_out_valid(PENetwork_56_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_56_io_to_pes_15_out_bits),
    .io_to_pes_15_sig_stat2trans(PENetwork_56_io_to_pes_15_sig_stat2trans),
    .io_to_pes_16_out_valid(PENetwork_56_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_56_io_to_pes_16_out_bits),
    .io_to_pes_16_sig_stat2trans(PENetwork_56_io_to_pes_16_sig_stat2trans),
    .io_to_pes_17_out_valid(PENetwork_56_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_56_io_to_pes_17_out_bits),
    .io_to_pes_17_sig_stat2trans(PENetwork_56_io_to_pes_17_sig_stat2trans),
    .io_to_pes_18_out_valid(PENetwork_56_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_56_io_to_pes_18_out_bits),
    .io_to_pes_18_sig_stat2trans(PENetwork_56_io_to_pes_18_sig_stat2trans),
    .io_to_pes_19_out_valid(PENetwork_56_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_56_io_to_pes_19_out_bits),
    .io_to_pes_19_sig_stat2trans(PENetwork_56_io_to_pes_19_sig_stat2trans),
    .io_to_pes_20_out_valid(PENetwork_56_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_56_io_to_pes_20_out_bits),
    .io_to_pes_20_sig_stat2trans(PENetwork_56_io_to_pes_20_sig_stat2trans),
    .io_to_pes_21_out_valid(PENetwork_56_io_to_pes_21_out_valid),
    .io_to_pes_21_out_bits(PENetwork_56_io_to_pes_21_out_bits),
    .io_to_pes_21_sig_stat2trans(PENetwork_56_io_to_pes_21_sig_stat2trans),
    .io_to_mem_valid(PENetwork_56_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_56_io_to_mem_bits),
    .io_sig_stat2trans(PENetwork_56_io_sig_stat2trans)
  );
  PENetwork_52 PENetwork_57 ( // @[pe.scala 229:13]
    .clock(PENetwork_57_clock),
    .reset(PENetwork_57_reset),
    .io_to_pes_0_out_valid(PENetwork_57_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_57_io_to_pes_0_out_bits),
    .io_to_pes_0_sig_stat2trans(PENetwork_57_io_to_pes_0_sig_stat2trans),
    .io_to_pes_1_out_valid(PENetwork_57_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_57_io_to_pes_1_out_bits),
    .io_to_pes_1_sig_stat2trans(PENetwork_57_io_to_pes_1_sig_stat2trans),
    .io_to_pes_2_out_valid(PENetwork_57_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_57_io_to_pes_2_out_bits),
    .io_to_pes_2_sig_stat2trans(PENetwork_57_io_to_pes_2_sig_stat2trans),
    .io_to_pes_3_out_valid(PENetwork_57_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_57_io_to_pes_3_out_bits),
    .io_to_pes_3_sig_stat2trans(PENetwork_57_io_to_pes_3_sig_stat2trans),
    .io_to_pes_4_out_valid(PENetwork_57_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_57_io_to_pes_4_out_bits),
    .io_to_pes_4_sig_stat2trans(PENetwork_57_io_to_pes_4_sig_stat2trans),
    .io_to_pes_5_out_valid(PENetwork_57_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_57_io_to_pes_5_out_bits),
    .io_to_pes_5_sig_stat2trans(PENetwork_57_io_to_pes_5_sig_stat2trans),
    .io_to_pes_6_out_valid(PENetwork_57_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_57_io_to_pes_6_out_bits),
    .io_to_pes_6_sig_stat2trans(PENetwork_57_io_to_pes_6_sig_stat2trans),
    .io_to_pes_7_out_valid(PENetwork_57_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_57_io_to_pes_7_out_bits),
    .io_to_pes_7_sig_stat2trans(PENetwork_57_io_to_pes_7_sig_stat2trans),
    .io_to_pes_8_out_valid(PENetwork_57_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_57_io_to_pes_8_out_bits),
    .io_to_pes_8_sig_stat2trans(PENetwork_57_io_to_pes_8_sig_stat2trans),
    .io_to_pes_9_out_valid(PENetwork_57_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_57_io_to_pes_9_out_bits),
    .io_to_pes_9_sig_stat2trans(PENetwork_57_io_to_pes_9_sig_stat2trans),
    .io_to_pes_10_out_valid(PENetwork_57_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_57_io_to_pes_10_out_bits),
    .io_to_pes_10_sig_stat2trans(PENetwork_57_io_to_pes_10_sig_stat2trans),
    .io_to_pes_11_out_valid(PENetwork_57_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_57_io_to_pes_11_out_bits),
    .io_to_pes_11_sig_stat2trans(PENetwork_57_io_to_pes_11_sig_stat2trans),
    .io_to_pes_12_out_valid(PENetwork_57_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_57_io_to_pes_12_out_bits),
    .io_to_pes_12_sig_stat2trans(PENetwork_57_io_to_pes_12_sig_stat2trans),
    .io_to_pes_13_out_valid(PENetwork_57_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_57_io_to_pes_13_out_bits),
    .io_to_pes_13_sig_stat2trans(PENetwork_57_io_to_pes_13_sig_stat2trans),
    .io_to_pes_14_out_valid(PENetwork_57_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_57_io_to_pes_14_out_bits),
    .io_to_pes_14_sig_stat2trans(PENetwork_57_io_to_pes_14_sig_stat2trans),
    .io_to_pes_15_out_valid(PENetwork_57_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_57_io_to_pes_15_out_bits),
    .io_to_pes_15_sig_stat2trans(PENetwork_57_io_to_pes_15_sig_stat2trans),
    .io_to_pes_16_out_valid(PENetwork_57_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_57_io_to_pes_16_out_bits),
    .io_to_pes_16_sig_stat2trans(PENetwork_57_io_to_pes_16_sig_stat2trans),
    .io_to_pes_17_out_valid(PENetwork_57_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_57_io_to_pes_17_out_bits),
    .io_to_pes_17_sig_stat2trans(PENetwork_57_io_to_pes_17_sig_stat2trans),
    .io_to_pes_18_out_valid(PENetwork_57_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_57_io_to_pes_18_out_bits),
    .io_to_pes_18_sig_stat2trans(PENetwork_57_io_to_pes_18_sig_stat2trans),
    .io_to_pes_19_out_valid(PENetwork_57_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_57_io_to_pes_19_out_bits),
    .io_to_pes_19_sig_stat2trans(PENetwork_57_io_to_pes_19_sig_stat2trans),
    .io_to_pes_20_out_valid(PENetwork_57_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_57_io_to_pes_20_out_bits),
    .io_to_pes_20_sig_stat2trans(PENetwork_57_io_to_pes_20_sig_stat2trans),
    .io_to_pes_21_out_valid(PENetwork_57_io_to_pes_21_out_valid),
    .io_to_pes_21_out_bits(PENetwork_57_io_to_pes_21_out_bits),
    .io_to_pes_21_sig_stat2trans(PENetwork_57_io_to_pes_21_sig_stat2trans),
    .io_to_mem_valid(PENetwork_57_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_57_io_to_mem_bits),
    .io_sig_stat2trans(PENetwork_57_io_sig_stat2trans)
  );
  PENetwork_52 PENetwork_58 ( // @[pe.scala 229:13]
    .clock(PENetwork_58_clock),
    .reset(PENetwork_58_reset),
    .io_to_pes_0_out_valid(PENetwork_58_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_58_io_to_pes_0_out_bits),
    .io_to_pes_0_sig_stat2trans(PENetwork_58_io_to_pes_0_sig_stat2trans),
    .io_to_pes_1_out_valid(PENetwork_58_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_58_io_to_pes_1_out_bits),
    .io_to_pes_1_sig_stat2trans(PENetwork_58_io_to_pes_1_sig_stat2trans),
    .io_to_pes_2_out_valid(PENetwork_58_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_58_io_to_pes_2_out_bits),
    .io_to_pes_2_sig_stat2trans(PENetwork_58_io_to_pes_2_sig_stat2trans),
    .io_to_pes_3_out_valid(PENetwork_58_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_58_io_to_pes_3_out_bits),
    .io_to_pes_3_sig_stat2trans(PENetwork_58_io_to_pes_3_sig_stat2trans),
    .io_to_pes_4_out_valid(PENetwork_58_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_58_io_to_pes_4_out_bits),
    .io_to_pes_4_sig_stat2trans(PENetwork_58_io_to_pes_4_sig_stat2trans),
    .io_to_pes_5_out_valid(PENetwork_58_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_58_io_to_pes_5_out_bits),
    .io_to_pes_5_sig_stat2trans(PENetwork_58_io_to_pes_5_sig_stat2trans),
    .io_to_pes_6_out_valid(PENetwork_58_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_58_io_to_pes_6_out_bits),
    .io_to_pes_6_sig_stat2trans(PENetwork_58_io_to_pes_6_sig_stat2trans),
    .io_to_pes_7_out_valid(PENetwork_58_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_58_io_to_pes_7_out_bits),
    .io_to_pes_7_sig_stat2trans(PENetwork_58_io_to_pes_7_sig_stat2trans),
    .io_to_pes_8_out_valid(PENetwork_58_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_58_io_to_pes_8_out_bits),
    .io_to_pes_8_sig_stat2trans(PENetwork_58_io_to_pes_8_sig_stat2trans),
    .io_to_pes_9_out_valid(PENetwork_58_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_58_io_to_pes_9_out_bits),
    .io_to_pes_9_sig_stat2trans(PENetwork_58_io_to_pes_9_sig_stat2trans),
    .io_to_pes_10_out_valid(PENetwork_58_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_58_io_to_pes_10_out_bits),
    .io_to_pes_10_sig_stat2trans(PENetwork_58_io_to_pes_10_sig_stat2trans),
    .io_to_pes_11_out_valid(PENetwork_58_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_58_io_to_pes_11_out_bits),
    .io_to_pes_11_sig_stat2trans(PENetwork_58_io_to_pes_11_sig_stat2trans),
    .io_to_pes_12_out_valid(PENetwork_58_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_58_io_to_pes_12_out_bits),
    .io_to_pes_12_sig_stat2trans(PENetwork_58_io_to_pes_12_sig_stat2trans),
    .io_to_pes_13_out_valid(PENetwork_58_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_58_io_to_pes_13_out_bits),
    .io_to_pes_13_sig_stat2trans(PENetwork_58_io_to_pes_13_sig_stat2trans),
    .io_to_pes_14_out_valid(PENetwork_58_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_58_io_to_pes_14_out_bits),
    .io_to_pes_14_sig_stat2trans(PENetwork_58_io_to_pes_14_sig_stat2trans),
    .io_to_pes_15_out_valid(PENetwork_58_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_58_io_to_pes_15_out_bits),
    .io_to_pes_15_sig_stat2trans(PENetwork_58_io_to_pes_15_sig_stat2trans),
    .io_to_pes_16_out_valid(PENetwork_58_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_58_io_to_pes_16_out_bits),
    .io_to_pes_16_sig_stat2trans(PENetwork_58_io_to_pes_16_sig_stat2trans),
    .io_to_pes_17_out_valid(PENetwork_58_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_58_io_to_pes_17_out_bits),
    .io_to_pes_17_sig_stat2trans(PENetwork_58_io_to_pes_17_sig_stat2trans),
    .io_to_pes_18_out_valid(PENetwork_58_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_58_io_to_pes_18_out_bits),
    .io_to_pes_18_sig_stat2trans(PENetwork_58_io_to_pes_18_sig_stat2trans),
    .io_to_pes_19_out_valid(PENetwork_58_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_58_io_to_pes_19_out_bits),
    .io_to_pes_19_sig_stat2trans(PENetwork_58_io_to_pes_19_sig_stat2trans),
    .io_to_pes_20_out_valid(PENetwork_58_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_58_io_to_pes_20_out_bits),
    .io_to_pes_20_sig_stat2trans(PENetwork_58_io_to_pes_20_sig_stat2trans),
    .io_to_pes_21_out_valid(PENetwork_58_io_to_pes_21_out_valid),
    .io_to_pes_21_out_bits(PENetwork_58_io_to_pes_21_out_bits),
    .io_to_pes_21_sig_stat2trans(PENetwork_58_io_to_pes_21_sig_stat2trans),
    .io_to_mem_valid(PENetwork_58_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_58_io_to_mem_bits),
    .io_sig_stat2trans(PENetwork_58_io_sig_stat2trans)
  );
  PENetwork_52 PENetwork_59 ( // @[pe.scala 229:13]
    .clock(PENetwork_59_clock),
    .reset(PENetwork_59_reset),
    .io_to_pes_0_out_valid(PENetwork_59_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_59_io_to_pes_0_out_bits),
    .io_to_pes_0_sig_stat2trans(PENetwork_59_io_to_pes_0_sig_stat2trans),
    .io_to_pes_1_out_valid(PENetwork_59_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_59_io_to_pes_1_out_bits),
    .io_to_pes_1_sig_stat2trans(PENetwork_59_io_to_pes_1_sig_stat2trans),
    .io_to_pes_2_out_valid(PENetwork_59_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_59_io_to_pes_2_out_bits),
    .io_to_pes_2_sig_stat2trans(PENetwork_59_io_to_pes_2_sig_stat2trans),
    .io_to_pes_3_out_valid(PENetwork_59_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_59_io_to_pes_3_out_bits),
    .io_to_pes_3_sig_stat2trans(PENetwork_59_io_to_pes_3_sig_stat2trans),
    .io_to_pes_4_out_valid(PENetwork_59_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_59_io_to_pes_4_out_bits),
    .io_to_pes_4_sig_stat2trans(PENetwork_59_io_to_pes_4_sig_stat2trans),
    .io_to_pes_5_out_valid(PENetwork_59_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_59_io_to_pes_5_out_bits),
    .io_to_pes_5_sig_stat2trans(PENetwork_59_io_to_pes_5_sig_stat2trans),
    .io_to_pes_6_out_valid(PENetwork_59_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_59_io_to_pes_6_out_bits),
    .io_to_pes_6_sig_stat2trans(PENetwork_59_io_to_pes_6_sig_stat2trans),
    .io_to_pes_7_out_valid(PENetwork_59_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_59_io_to_pes_7_out_bits),
    .io_to_pes_7_sig_stat2trans(PENetwork_59_io_to_pes_7_sig_stat2trans),
    .io_to_pes_8_out_valid(PENetwork_59_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_59_io_to_pes_8_out_bits),
    .io_to_pes_8_sig_stat2trans(PENetwork_59_io_to_pes_8_sig_stat2trans),
    .io_to_pes_9_out_valid(PENetwork_59_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_59_io_to_pes_9_out_bits),
    .io_to_pes_9_sig_stat2trans(PENetwork_59_io_to_pes_9_sig_stat2trans),
    .io_to_pes_10_out_valid(PENetwork_59_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_59_io_to_pes_10_out_bits),
    .io_to_pes_10_sig_stat2trans(PENetwork_59_io_to_pes_10_sig_stat2trans),
    .io_to_pes_11_out_valid(PENetwork_59_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_59_io_to_pes_11_out_bits),
    .io_to_pes_11_sig_stat2trans(PENetwork_59_io_to_pes_11_sig_stat2trans),
    .io_to_pes_12_out_valid(PENetwork_59_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_59_io_to_pes_12_out_bits),
    .io_to_pes_12_sig_stat2trans(PENetwork_59_io_to_pes_12_sig_stat2trans),
    .io_to_pes_13_out_valid(PENetwork_59_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_59_io_to_pes_13_out_bits),
    .io_to_pes_13_sig_stat2trans(PENetwork_59_io_to_pes_13_sig_stat2trans),
    .io_to_pes_14_out_valid(PENetwork_59_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_59_io_to_pes_14_out_bits),
    .io_to_pes_14_sig_stat2trans(PENetwork_59_io_to_pes_14_sig_stat2trans),
    .io_to_pes_15_out_valid(PENetwork_59_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_59_io_to_pes_15_out_bits),
    .io_to_pes_15_sig_stat2trans(PENetwork_59_io_to_pes_15_sig_stat2trans),
    .io_to_pes_16_out_valid(PENetwork_59_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_59_io_to_pes_16_out_bits),
    .io_to_pes_16_sig_stat2trans(PENetwork_59_io_to_pes_16_sig_stat2trans),
    .io_to_pes_17_out_valid(PENetwork_59_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_59_io_to_pes_17_out_bits),
    .io_to_pes_17_sig_stat2trans(PENetwork_59_io_to_pes_17_sig_stat2trans),
    .io_to_pes_18_out_valid(PENetwork_59_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_59_io_to_pes_18_out_bits),
    .io_to_pes_18_sig_stat2trans(PENetwork_59_io_to_pes_18_sig_stat2trans),
    .io_to_pes_19_out_valid(PENetwork_59_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_59_io_to_pes_19_out_bits),
    .io_to_pes_19_sig_stat2trans(PENetwork_59_io_to_pes_19_sig_stat2trans),
    .io_to_pes_20_out_valid(PENetwork_59_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_59_io_to_pes_20_out_bits),
    .io_to_pes_20_sig_stat2trans(PENetwork_59_io_to_pes_20_sig_stat2trans),
    .io_to_pes_21_out_valid(PENetwork_59_io_to_pes_21_out_valid),
    .io_to_pes_21_out_bits(PENetwork_59_io_to_pes_21_out_bits),
    .io_to_pes_21_sig_stat2trans(PENetwork_59_io_to_pes_21_sig_stat2trans),
    .io_to_mem_valid(PENetwork_59_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_59_io_to_mem_bits),
    .io_sig_stat2trans(PENetwork_59_io_sig_stat2trans)
  );
  PENetwork_52 PENetwork_60 ( // @[pe.scala 229:13]
    .clock(PENetwork_60_clock),
    .reset(PENetwork_60_reset),
    .io_to_pes_0_out_valid(PENetwork_60_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_60_io_to_pes_0_out_bits),
    .io_to_pes_0_sig_stat2trans(PENetwork_60_io_to_pes_0_sig_stat2trans),
    .io_to_pes_1_out_valid(PENetwork_60_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_60_io_to_pes_1_out_bits),
    .io_to_pes_1_sig_stat2trans(PENetwork_60_io_to_pes_1_sig_stat2trans),
    .io_to_pes_2_out_valid(PENetwork_60_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_60_io_to_pes_2_out_bits),
    .io_to_pes_2_sig_stat2trans(PENetwork_60_io_to_pes_2_sig_stat2trans),
    .io_to_pes_3_out_valid(PENetwork_60_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_60_io_to_pes_3_out_bits),
    .io_to_pes_3_sig_stat2trans(PENetwork_60_io_to_pes_3_sig_stat2trans),
    .io_to_pes_4_out_valid(PENetwork_60_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_60_io_to_pes_4_out_bits),
    .io_to_pes_4_sig_stat2trans(PENetwork_60_io_to_pes_4_sig_stat2trans),
    .io_to_pes_5_out_valid(PENetwork_60_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_60_io_to_pes_5_out_bits),
    .io_to_pes_5_sig_stat2trans(PENetwork_60_io_to_pes_5_sig_stat2trans),
    .io_to_pes_6_out_valid(PENetwork_60_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_60_io_to_pes_6_out_bits),
    .io_to_pes_6_sig_stat2trans(PENetwork_60_io_to_pes_6_sig_stat2trans),
    .io_to_pes_7_out_valid(PENetwork_60_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_60_io_to_pes_7_out_bits),
    .io_to_pes_7_sig_stat2trans(PENetwork_60_io_to_pes_7_sig_stat2trans),
    .io_to_pes_8_out_valid(PENetwork_60_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_60_io_to_pes_8_out_bits),
    .io_to_pes_8_sig_stat2trans(PENetwork_60_io_to_pes_8_sig_stat2trans),
    .io_to_pes_9_out_valid(PENetwork_60_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_60_io_to_pes_9_out_bits),
    .io_to_pes_9_sig_stat2trans(PENetwork_60_io_to_pes_9_sig_stat2trans),
    .io_to_pes_10_out_valid(PENetwork_60_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_60_io_to_pes_10_out_bits),
    .io_to_pes_10_sig_stat2trans(PENetwork_60_io_to_pes_10_sig_stat2trans),
    .io_to_pes_11_out_valid(PENetwork_60_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_60_io_to_pes_11_out_bits),
    .io_to_pes_11_sig_stat2trans(PENetwork_60_io_to_pes_11_sig_stat2trans),
    .io_to_pes_12_out_valid(PENetwork_60_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_60_io_to_pes_12_out_bits),
    .io_to_pes_12_sig_stat2trans(PENetwork_60_io_to_pes_12_sig_stat2trans),
    .io_to_pes_13_out_valid(PENetwork_60_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_60_io_to_pes_13_out_bits),
    .io_to_pes_13_sig_stat2trans(PENetwork_60_io_to_pes_13_sig_stat2trans),
    .io_to_pes_14_out_valid(PENetwork_60_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_60_io_to_pes_14_out_bits),
    .io_to_pes_14_sig_stat2trans(PENetwork_60_io_to_pes_14_sig_stat2trans),
    .io_to_pes_15_out_valid(PENetwork_60_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_60_io_to_pes_15_out_bits),
    .io_to_pes_15_sig_stat2trans(PENetwork_60_io_to_pes_15_sig_stat2trans),
    .io_to_pes_16_out_valid(PENetwork_60_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_60_io_to_pes_16_out_bits),
    .io_to_pes_16_sig_stat2trans(PENetwork_60_io_to_pes_16_sig_stat2trans),
    .io_to_pes_17_out_valid(PENetwork_60_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_60_io_to_pes_17_out_bits),
    .io_to_pes_17_sig_stat2trans(PENetwork_60_io_to_pes_17_sig_stat2trans),
    .io_to_pes_18_out_valid(PENetwork_60_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_60_io_to_pes_18_out_bits),
    .io_to_pes_18_sig_stat2trans(PENetwork_60_io_to_pes_18_sig_stat2trans),
    .io_to_pes_19_out_valid(PENetwork_60_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_60_io_to_pes_19_out_bits),
    .io_to_pes_19_sig_stat2trans(PENetwork_60_io_to_pes_19_sig_stat2trans),
    .io_to_pes_20_out_valid(PENetwork_60_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_60_io_to_pes_20_out_bits),
    .io_to_pes_20_sig_stat2trans(PENetwork_60_io_to_pes_20_sig_stat2trans),
    .io_to_pes_21_out_valid(PENetwork_60_io_to_pes_21_out_valid),
    .io_to_pes_21_out_bits(PENetwork_60_io_to_pes_21_out_bits),
    .io_to_pes_21_sig_stat2trans(PENetwork_60_io_to_pes_21_sig_stat2trans),
    .io_to_mem_valid(PENetwork_60_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_60_io_to_mem_bits),
    .io_sig_stat2trans(PENetwork_60_io_sig_stat2trans)
  );
  PENetwork_52 PENetwork_61 ( // @[pe.scala 229:13]
    .clock(PENetwork_61_clock),
    .reset(PENetwork_61_reset),
    .io_to_pes_0_out_valid(PENetwork_61_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_61_io_to_pes_0_out_bits),
    .io_to_pes_0_sig_stat2trans(PENetwork_61_io_to_pes_0_sig_stat2trans),
    .io_to_pes_1_out_valid(PENetwork_61_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_61_io_to_pes_1_out_bits),
    .io_to_pes_1_sig_stat2trans(PENetwork_61_io_to_pes_1_sig_stat2trans),
    .io_to_pes_2_out_valid(PENetwork_61_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_61_io_to_pes_2_out_bits),
    .io_to_pes_2_sig_stat2trans(PENetwork_61_io_to_pes_2_sig_stat2trans),
    .io_to_pes_3_out_valid(PENetwork_61_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_61_io_to_pes_3_out_bits),
    .io_to_pes_3_sig_stat2trans(PENetwork_61_io_to_pes_3_sig_stat2trans),
    .io_to_pes_4_out_valid(PENetwork_61_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_61_io_to_pes_4_out_bits),
    .io_to_pes_4_sig_stat2trans(PENetwork_61_io_to_pes_4_sig_stat2trans),
    .io_to_pes_5_out_valid(PENetwork_61_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_61_io_to_pes_5_out_bits),
    .io_to_pes_5_sig_stat2trans(PENetwork_61_io_to_pes_5_sig_stat2trans),
    .io_to_pes_6_out_valid(PENetwork_61_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_61_io_to_pes_6_out_bits),
    .io_to_pes_6_sig_stat2trans(PENetwork_61_io_to_pes_6_sig_stat2trans),
    .io_to_pes_7_out_valid(PENetwork_61_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_61_io_to_pes_7_out_bits),
    .io_to_pes_7_sig_stat2trans(PENetwork_61_io_to_pes_7_sig_stat2trans),
    .io_to_pes_8_out_valid(PENetwork_61_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_61_io_to_pes_8_out_bits),
    .io_to_pes_8_sig_stat2trans(PENetwork_61_io_to_pes_8_sig_stat2trans),
    .io_to_pes_9_out_valid(PENetwork_61_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_61_io_to_pes_9_out_bits),
    .io_to_pes_9_sig_stat2trans(PENetwork_61_io_to_pes_9_sig_stat2trans),
    .io_to_pes_10_out_valid(PENetwork_61_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_61_io_to_pes_10_out_bits),
    .io_to_pes_10_sig_stat2trans(PENetwork_61_io_to_pes_10_sig_stat2trans),
    .io_to_pes_11_out_valid(PENetwork_61_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_61_io_to_pes_11_out_bits),
    .io_to_pes_11_sig_stat2trans(PENetwork_61_io_to_pes_11_sig_stat2trans),
    .io_to_pes_12_out_valid(PENetwork_61_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_61_io_to_pes_12_out_bits),
    .io_to_pes_12_sig_stat2trans(PENetwork_61_io_to_pes_12_sig_stat2trans),
    .io_to_pes_13_out_valid(PENetwork_61_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_61_io_to_pes_13_out_bits),
    .io_to_pes_13_sig_stat2trans(PENetwork_61_io_to_pes_13_sig_stat2trans),
    .io_to_pes_14_out_valid(PENetwork_61_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_61_io_to_pes_14_out_bits),
    .io_to_pes_14_sig_stat2trans(PENetwork_61_io_to_pes_14_sig_stat2trans),
    .io_to_pes_15_out_valid(PENetwork_61_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_61_io_to_pes_15_out_bits),
    .io_to_pes_15_sig_stat2trans(PENetwork_61_io_to_pes_15_sig_stat2trans),
    .io_to_pes_16_out_valid(PENetwork_61_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_61_io_to_pes_16_out_bits),
    .io_to_pes_16_sig_stat2trans(PENetwork_61_io_to_pes_16_sig_stat2trans),
    .io_to_pes_17_out_valid(PENetwork_61_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_61_io_to_pes_17_out_bits),
    .io_to_pes_17_sig_stat2trans(PENetwork_61_io_to_pes_17_sig_stat2trans),
    .io_to_pes_18_out_valid(PENetwork_61_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_61_io_to_pes_18_out_bits),
    .io_to_pes_18_sig_stat2trans(PENetwork_61_io_to_pes_18_sig_stat2trans),
    .io_to_pes_19_out_valid(PENetwork_61_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_61_io_to_pes_19_out_bits),
    .io_to_pes_19_sig_stat2trans(PENetwork_61_io_to_pes_19_sig_stat2trans),
    .io_to_pes_20_out_valid(PENetwork_61_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_61_io_to_pes_20_out_bits),
    .io_to_pes_20_sig_stat2trans(PENetwork_61_io_to_pes_20_sig_stat2trans),
    .io_to_pes_21_out_valid(PENetwork_61_io_to_pes_21_out_valid),
    .io_to_pes_21_out_bits(PENetwork_61_io_to_pes_21_out_bits),
    .io_to_pes_21_sig_stat2trans(PENetwork_61_io_to_pes_21_sig_stat2trans),
    .io_to_mem_valid(PENetwork_61_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_61_io_to_mem_bits),
    .io_sig_stat2trans(PENetwork_61_io_sig_stat2trans)
  );
  PENetwork_52 PENetwork_62 ( // @[pe.scala 229:13]
    .clock(PENetwork_62_clock),
    .reset(PENetwork_62_reset),
    .io_to_pes_0_out_valid(PENetwork_62_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_62_io_to_pes_0_out_bits),
    .io_to_pes_0_sig_stat2trans(PENetwork_62_io_to_pes_0_sig_stat2trans),
    .io_to_pes_1_out_valid(PENetwork_62_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_62_io_to_pes_1_out_bits),
    .io_to_pes_1_sig_stat2trans(PENetwork_62_io_to_pes_1_sig_stat2trans),
    .io_to_pes_2_out_valid(PENetwork_62_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_62_io_to_pes_2_out_bits),
    .io_to_pes_2_sig_stat2trans(PENetwork_62_io_to_pes_2_sig_stat2trans),
    .io_to_pes_3_out_valid(PENetwork_62_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_62_io_to_pes_3_out_bits),
    .io_to_pes_3_sig_stat2trans(PENetwork_62_io_to_pes_3_sig_stat2trans),
    .io_to_pes_4_out_valid(PENetwork_62_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_62_io_to_pes_4_out_bits),
    .io_to_pes_4_sig_stat2trans(PENetwork_62_io_to_pes_4_sig_stat2trans),
    .io_to_pes_5_out_valid(PENetwork_62_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_62_io_to_pes_5_out_bits),
    .io_to_pes_5_sig_stat2trans(PENetwork_62_io_to_pes_5_sig_stat2trans),
    .io_to_pes_6_out_valid(PENetwork_62_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_62_io_to_pes_6_out_bits),
    .io_to_pes_6_sig_stat2trans(PENetwork_62_io_to_pes_6_sig_stat2trans),
    .io_to_pes_7_out_valid(PENetwork_62_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_62_io_to_pes_7_out_bits),
    .io_to_pes_7_sig_stat2trans(PENetwork_62_io_to_pes_7_sig_stat2trans),
    .io_to_pes_8_out_valid(PENetwork_62_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_62_io_to_pes_8_out_bits),
    .io_to_pes_8_sig_stat2trans(PENetwork_62_io_to_pes_8_sig_stat2trans),
    .io_to_pes_9_out_valid(PENetwork_62_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_62_io_to_pes_9_out_bits),
    .io_to_pes_9_sig_stat2trans(PENetwork_62_io_to_pes_9_sig_stat2trans),
    .io_to_pes_10_out_valid(PENetwork_62_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_62_io_to_pes_10_out_bits),
    .io_to_pes_10_sig_stat2trans(PENetwork_62_io_to_pes_10_sig_stat2trans),
    .io_to_pes_11_out_valid(PENetwork_62_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_62_io_to_pes_11_out_bits),
    .io_to_pes_11_sig_stat2trans(PENetwork_62_io_to_pes_11_sig_stat2trans),
    .io_to_pes_12_out_valid(PENetwork_62_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_62_io_to_pes_12_out_bits),
    .io_to_pes_12_sig_stat2trans(PENetwork_62_io_to_pes_12_sig_stat2trans),
    .io_to_pes_13_out_valid(PENetwork_62_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_62_io_to_pes_13_out_bits),
    .io_to_pes_13_sig_stat2trans(PENetwork_62_io_to_pes_13_sig_stat2trans),
    .io_to_pes_14_out_valid(PENetwork_62_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_62_io_to_pes_14_out_bits),
    .io_to_pes_14_sig_stat2trans(PENetwork_62_io_to_pes_14_sig_stat2trans),
    .io_to_pes_15_out_valid(PENetwork_62_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_62_io_to_pes_15_out_bits),
    .io_to_pes_15_sig_stat2trans(PENetwork_62_io_to_pes_15_sig_stat2trans),
    .io_to_pes_16_out_valid(PENetwork_62_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_62_io_to_pes_16_out_bits),
    .io_to_pes_16_sig_stat2trans(PENetwork_62_io_to_pes_16_sig_stat2trans),
    .io_to_pes_17_out_valid(PENetwork_62_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_62_io_to_pes_17_out_bits),
    .io_to_pes_17_sig_stat2trans(PENetwork_62_io_to_pes_17_sig_stat2trans),
    .io_to_pes_18_out_valid(PENetwork_62_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_62_io_to_pes_18_out_bits),
    .io_to_pes_18_sig_stat2trans(PENetwork_62_io_to_pes_18_sig_stat2trans),
    .io_to_pes_19_out_valid(PENetwork_62_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_62_io_to_pes_19_out_bits),
    .io_to_pes_19_sig_stat2trans(PENetwork_62_io_to_pes_19_sig_stat2trans),
    .io_to_pes_20_out_valid(PENetwork_62_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_62_io_to_pes_20_out_bits),
    .io_to_pes_20_sig_stat2trans(PENetwork_62_io_to_pes_20_sig_stat2trans),
    .io_to_pes_21_out_valid(PENetwork_62_io_to_pes_21_out_valid),
    .io_to_pes_21_out_bits(PENetwork_62_io_to_pes_21_out_bits),
    .io_to_pes_21_sig_stat2trans(PENetwork_62_io_to_pes_21_sig_stat2trans),
    .io_to_mem_valid(PENetwork_62_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_62_io_to_mem_bits),
    .io_sig_stat2trans(PENetwork_62_io_sig_stat2trans)
  );
  PENetwork_52 PENetwork_63 ( // @[pe.scala 229:13]
    .clock(PENetwork_63_clock),
    .reset(PENetwork_63_reset),
    .io_to_pes_0_out_valid(PENetwork_63_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_63_io_to_pes_0_out_bits),
    .io_to_pes_0_sig_stat2trans(PENetwork_63_io_to_pes_0_sig_stat2trans),
    .io_to_pes_1_out_valid(PENetwork_63_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_63_io_to_pes_1_out_bits),
    .io_to_pes_1_sig_stat2trans(PENetwork_63_io_to_pes_1_sig_stat2trans),
    .io_to_pes_2_out_valid(PENetwork_63_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_63_io_to_pes_2_out_bits),
    .io_to_pes_2_sig_stat2trans(PENetwork_63_io_to_pes_2_sig_stat2trans),
    .io_to_pes_3_out_valid(PENetwork_63_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_63_io_to_pes_3_out_bits),
    .io_to_pes_3_sig_stat2trans(PENetwork_63_io_to_pes_3_sig_stat2trans),
    .io_to_pes_4_out_valid(PENetwork_63_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_63_io_to_pes_4_out_bits),
    .io_to_pes_4_sig_stat2trans(PENetwork_63_io_to_pes_4_sig_stat2trans),
    .io_to_pes_5_out_valid(PENetwork_63_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_63_io_to_pes_5_out_bits),
    .io_to_pes_5_sig_stat2trans(PENetwork_63_io_to_pes_5_sig_stat2trans),
    .io_to_pes_6_out_valid(PENetwork_63_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_63_io_to_pes_6_out_bits),
    .io_to_pes_6_sig_stat2trans(PENetwork_63_io_to_pes_6_sig_stat2trans),
    .io_to_pes_7_out_valid(PENetwork_63_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_63_io_to_pes_7_out_bits),
    .io_to_pes_7_sig_stat2trans(PENetwork_63_io_to_pes_7_sig_stat2trans),
    .io_to_pes_8_out_valid(PENetwork_63_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_63_io_to_pes_8_out_bits),
    .io_to_pes_8_sig_stat2trans(PENetwork_63_io_to_pes_8_sig_stat2trans),
    .io_to_pes_9_out_valid(PENetwork_63_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_63_io_to_pes_9_out_bits),
    .io_to_pes_9_sig_stat2trans(PENetwork_63_io_to_pes_9_sig_stat2trans),
    .io_to_pes_10_out_valid(PENetwork_63_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_63_io_to_pes_10_out_bits),
    .io_to_pes_10_sig_stat2trans(PENetwork_63_io_to_pes_10_sig_stat2trans),
    .io_to_pes_11_out_valid(PENetwork_63_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_63_io_to_pes_11_out_bits),
    .io_to_pes_11_sig_stat2trans(PENetwork_63_io_to_pes_11_sig_stat2trans),
    .io_to_pes_12_out_valid(PENetwork_63_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_63_io_to_pes_12_out_bits),
    .io_to_pes_12_sig_stat2trans(PENetwork_63_io_to_pes_12_sig_stat2trans),
    .io_to_pes_13_out_valid(PENetwork_63_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_63_io_to_pes_13_out_bits),
    .io_to_pes_13_sig_stat2trans(PENetwork_63_io_to_pes_13_sig_stat2trans),
    .io_to_pes_14_out_valid(PENetwork_63_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_63_io_to_pes_14_out_bits),
    .io_to_pes_14_sig_stat2trans(PENetwork_63_io_to_pes_14_sig_stat2trans),
    .io_to_pes_15_out_valid(PENetwork_63_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_63_io_to_pes_15_out_bits),
    .io_to_pes_15_sig_stat2trans(PENetwork_63_io_to_pes_15_sig_stat2trans),
    .io_to_pes_16_out_valid(PENetwork_63_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_63_io_to_pes_16_out_bits),
    .io_to_pes_16_sig_stat2trans(PENetwork_63_io_to_pes_16_sig_stat2trans),
    .io_to_pes_17_out_valid(PENetwork_63_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_63_io_to_pes_17_out_bits),
    .io_to_pes_17_sig_stat2trans(PENetwork_63_io_to_pes_17_sig_stat2trans),
    .io_to_pes_18_out_valid(PENetwork_63_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_63_io_to_pes_18_out_bits),
    .io_to_pes_18_sig_stat2trans(PENetwork_63_io_to_pes_18_sig_stat2trans),
    .io_to_pes_19_out_valid(PENetwork_63_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_63_io_to_pes_19_out_bits),
    .io_to_pes_19_sig_stat2trans(PENetwork_63_io_to_pes_19_sig_stat2trans),
    .io_to_pes_20_out_valid(PENetwork_63_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_63_io_to_pes_20_out_bits),
    .io_to_pes_20_sig_stat2trans(PENetwork_63_io_to_pes_20_sig_stat2trans),
    .io_to_pes_21_out_valid(PENetwork_63_io_to_pes_21_out_valid),
    .io_to_pes_21_out_bits(PENetwork_63_io_to_pes_21_out_bits),
    .io_to_pes_21_sig_stat2trans(PENetwork_63_io_to_pes_21_sig_stat2trans),
    .io_to_mem_valid(PENetwork_63_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_63_io_to_mem_bits),
    .io_sig_stat2trans(PENetwork_63_io_sig_stat2trans)
  );
  PENetwork_52 PENetwork_64 ( // @[pe.scala 229:13]
    .clock(PENetwork_64_clock),
    .reset(PENetwork_64_reset),
    .io_to_pes_0_out_valid(PENetwork_64_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_64_io_to_pes_0_out_bits),
    .io_to_pes_0_sig_stat2trans(PENetwork_64_io_to_pes_0_sig_stat2trans),
    .io_to_pes_1_out_valid(PENetwork_64_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_64_io_to_pes_1_out_bits),
    .io_to_pes_1_sig_stat2trans(PENetwork_64_io_to_pes_1_sig_stat2trans),
    .io_to_pes_2_out_valid(PENetwork_64_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_64_io_to_pes_2_out_bits),
    .io_to_pes_2_sig_stat2trans(PENetwork_64_io_to_pes_2_sig_stat2trans),
    .io_to_pes_3_out_valid(PENetwork_64_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_64_io_to_pes_3_out_bits),
    .io_to_pes_3_sig_stat2trans(PENetwork_64_io_to_pes_3_sig_stat2trans),
    .io_to_pes_4_out_valid(PENetwork_64_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_64_io_to_pes_4_out_bits),
    .io_to_pes_4_sig_stat2trans(PENetwork_64_io_to_pes_4_sig_stat2trans),
    .io_to_pes_5_out_valid(PENetwork_64_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_64_io_to_pes_5_out_bits),
    .io_to_pes_5_sig_stat2trans(PENetwork_64_io_to_pes_5_sig_stat2trans),
    .io_to_pes_6_out_valid(PENetwork_64_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_64_io_to_pes_6_out_bits),
    .io_to_pes_6_sig_stat2trans(PENetwork_64_io_to_pes_6_sig_stat2trans),
    .io_to_pes_7_out_valid(PENetwork_64_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_64_io_to_pes_7_out_bits),
    .io_to_pes_7_sig_stat2trans(PENetwork_64_io_to_pes_7_sig_stat2trans),
    .io_to_pes_8_out_valid(PENetwork_64_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_64_io_to_pes_8_out_bits),
    .io_to_pes_8_sig_stat2trans(PENetwork_64_io_to_pes_8_sig_stat2trans),
    .io_to_pes_9_out_valid(PENetwork_64_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_64_io_to_pes_9_out_bits),
    .io_to_pes_9_sig_stat2trans(PENetwork_64_io_to_pes_9_sig_stat2trans),
    .io_to_pes_10_out_valid(PENetwork_64_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_64_io_to_pes_10_out_bits),
    .io_to_pes_10_sig_stat2trans(PENetwork_64_io_to_pes_10_sig_stat2trans),
    .io_to_pes_11_out_valid(PENetwork_64_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_64_io_to_pes_11_out_bits),
    .io_to_pes_11_sig_stat2trans(PENetwork_64_io_to_pes_11_sig_stat2trans),
    .io_to_pes_12_out_valid(PENetwork_64_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_64_io_to_pes_12_out_bits),
    .io_to_pes_12_sig_stat2trans(PENetwork_64_io_to_pes_12_sig_stat2trans),
    .io_to_pes_13_out_valid(PENetwork_64_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_64_io_to_pes_13_out_bits),
    .io_to_pes_13_sig_stat2trans(PENetwork_64_io_to_pes_13_sig_stat2trans),
    .io_to_pes_14_out_valid(PENetwork_64_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_64_io_to_pes_14_out_bits),
    .io_to_pes_14_sig_stat2trans(PENetwork_64_io_to_pes_14_sig_stat2trans),
    .io_to_pes_15_out_valid(PENetwork_64_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_64_io_to_pes_15_out_bits),
    .io_to_pes_15_sig_stat2trans(PENetwork_64_io_to_pes_15_sig_stat2trans),
    .io_to_pes_16_out_valid(PENetwork_64_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_64_io_to_pes_16_out_bits),
    .io_to_pes_16_sig_stat2trans(PENetwork_64_io_to_pes_16_sig_stat2trans),
    .io_to_pes_17_out_valid(PENetwork_64_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_64_io_to_pes_17_out_bits),
    .io_to_pes_17_sig_stat2trans(PENetwork_64_io_to_pes_17_sig_stat2trans),
    .io_to_pes_18_out_valid(PENetwork_64_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_64_io_to_pes_18_out_bits),
    .io_to_pes_18_sig_stat2trans(PENetwork_64_io_to_pes_18_sig_stat2trans),
    .io_to_pes_19_out_valid(PENetwork_64_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_64_io_to_pes_19_out_bits),
    .io_to_pes_19_sig_stat2trans(PENetwork_64_io_to_pes_19_sig_stat2trans),
    .io_to_pes_20_out_valid(PENetwork_64_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_64_io_to_pes_20_out_bits),
    .io_to_pes_20_sig_stat2trans(PENetwork_64_io_to_pes_20_sig_stat2trans),
    .io_to_pes_21_out_valid(PENetwork_64_io_to_pes_21_out_valid),
    .io_to_pes_21_out_bits(PENetwork_64_io_to_pes_21_out_bits),
    .io_to_pes_21_sig_stat2trans(PENetwork_64_io_to_pes_21_sig_stat2trans),
    .io_to_mem_valid(PENetwork_64_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_64_io_to_mem_bits),
    .io_sig_stat2trans(PENetwork_64_io_sig_stat2trans)
  );
  PENetwork_52 PENetwork_65 ( // @[pe.scala 229:13]
    .clock(PENetwork_65_clock),
    .reset(PENetwork_65_reset),
    .io_to_pes_0_out_valid(PENetwork_65_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_65_io_to_pes_0_out_bits),
    .io_to_pes_0_sig_stat2trans(PENetwork_65_io_to_pes_0_sig_stat2trans),
    .io_to_pes_1_out_valid(PENetwork_65_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_65_io_to_pes_1_out_bits),
    .io_to_pes_1_sig_stat2trans(PENetwork_65_io_to_pes_1_sig_stat2trans),
    .io_to_pes_2_out_valid(PENetwork_65_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_65_io_to_pes_2_out_bits),
    .io_to_pes_2_sig_stat2trans(PENetwork_65_io_to_pes_2_sig_stat2trans),
    .io_to_pes_3_out_valid(PENetwork_65_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_65_io_to_pes_3_out_bits),
    .io_to_pes_3_sig_stat2trans(PENetwork_65_io_to_pes_3_sig_stat2trans),
    .io_to_pes_4_out_valid(PENetwork_65_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_65_io_to_pes_4_out_bits),
    .io_to_pes_4_sig_stat2trans(PENetwork_65_io_to_pes_4_sig_stat2trans),
    .io_to_pes_5_out_valid(PENetwork_65_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_65_io_to_pes_5_out_bits),
    .io_to_pes_5_sig_stat2trans(PENetwork_65_io_to_pes_5_sig_stat2trans),
    .io_to_pes_6_out_valid(PENetwork_65_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_65_io_to_pes_6_out_bits),
    .io_to_pes_6_sig_stat2trans(PENetwork_65_io_to_pes_6_sig_stat2trans),
    .io_to_pes_7_out_valid(PENetwork_65_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_65_io_to_pes_7_out_bits),
    .io_to_pes_7_sig_stat2trans(PENetwork_65_io_to_pes_7_sig_stat2trans),
    .io_to_pes_8_out_valid(PENetwork_65_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_65_io_to_pes_8_out_bits),
    .io_to_pes_8_sig_stat2trans(PENetwork_65_io_to_pes_8_sig_stat2trans),
    .io_to_pes_9_out_valid(PENetwork_65_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_65_io_to_pes_9_out_bits),
    .io_to_pes_9_sig_stat2trans(PENetwork_65_io_to_pes_9_sig_stat2trans),
    .io_to_pes_10_out_valid(PENetwork_65_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_65_io_to_pes_10_out_bits),
    .io_to_pes_10_sig_stat2trans(PENetwork_65_io_to_pes_10_sig_stat2trans),
    .io_to_pes_11_out_valid(PENetwork_65_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_65_io_to_pes_11_out_bits),
    .io_to_pes_11_sig_stat2trans(PENetwork_65_io_to_pes_11_sig_stat2trans),
    .io_to_pes_12_out_valid(PENetwork_65_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_65_io_to_pes_12_out_bits),
    .io_to_pes_12_sig_stat2trans(PENetwork_65_io_to_pes_12_sig_stat2trans),
    .io_to_pes_13_out_valid(PENetwork_65_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_65_io_to_pes_13_out_bits),
    .io_to_pes_13_sig_stat2trans(PENetwork_65_io_to_pes_13_sig_stat2trans),
    .io_to_pes_14_out_valid(PENetwork_65_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_65_io_to_pes_14_out_bits),
    .io_to_pes_14_sig_stat2trans(PENetwork_65_io_to_pes_14_sig_stat2trans),
    .io_to_pes_15_out_valid(PENetwork_65_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_65_io_to_pes_15_out_bits),
    .io_to_pes_15_sig_stat2trans(PENetwork_65_io_to_pes_15_sig_stat2trans),
    .io_to_pes_16_out_valid(PENetwork_65_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_65_io_to_pes_16_out_bits),
    .io_to_pes_16_sig_stat2trans(PENetwork_65_io_to_pes_16_sig_stat2trans),
    .io_to_pes_17_out_valid(PENetwork_65_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_65_io_to_pes_17_out_bits),
    .io_to_pes_17_sig_stat2trans(PENetwork_65_io_to_pes_17_sig_stat2trans),
    .io_to_pes_18_out_valid(PENetwork_65_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_65_io_to_pes_18_out_bits),
    .io_to_pes_18_sig_stat2trans(PENetwork_65_io_to_pes_18_sig_stat2trans),
    .io_to_pes_19_out_valid(PENetwork_65_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_65_io_to_pes_19_out_bits),
    .io_to_pes_19_sig_stat2trans(PENetwork_65_io_to_pes_19_sig_stat2trans),
    .io_to_pes_20_out_valid(PENetwork_65_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_65_io_to_pes_20_out_bits),
    .io_to_pes_20_sig_stat2trans(PENetwork_65_io_to_pes_20_sig_stat2trans),
    .io_to_pes_21_out_valid(PENetwork_65_io_to_pes_21_out_valid),
    .io_to_pes_21_out_bits(PENetwork_65_io_to_pes_21_out_bits),
    .io_to_pes_21_sig_stat2trans(PENetwork_65_io_to_pes_21_sig_stat2trans),
    .io_to_mem_valid(PENetwork_65_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_65_io_to_mem_bits),
    .io_sig_stat2trans(PENetwork_65_io_sig_stat2trans)
  );
  PENetwork_52 PENetwork_66 ( // @[pe.scala 229:13]
    .clock(PENetwork_66_clock),
    .reset(PENetwork_66_reset),
    .io_to_pes_0_out_valid(PENetwork_66_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_66_io_to_pes_0_out_bits),
    .io_to_pes_0_sig_stat2trans(PENetwork_66_io_to_pes_0_sig_stat2trans),
    .io_to_pes_1_out_valid(PENetwork_66_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_66_io_to_pes_1_out_bits),
    .io_to_pes_1_sig_stat2trans(PENetwork_66_io_to_pes_1_sig_stat2trans),
    .io_to_pes_2_out_valid(PENetwork_66_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_66_io_to_pes_2_out_bits),
    .io_to_pes_2_sig_stat2trans(PENetwork_66_io_to_pes_2_sig_stat2trans),
    .io_to_pes_3_out_valid(PENetwork_66_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_66_io_to_pes_3_out_bits),
    .io_to_pes_3_sig_stat2trans(PENetwork_66_io_to_pes_3_sig_stat2trans),
    .io_to_pes_4_out_valid(PENetwork_66_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_66_io_to_pes_4_out_bits),
    .io_to_pes_4_sig_stat2trans(PENetwork_66_io_to_pes_4_sig_stat2trans),
    .io_to_pes_5_out_valid(PENetwork_66_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_66_io_to_pes_5_out_bits),
    .io_to_pes_5_sig_stat2trans(PENetwork_66_io_to_pes_5_sig_stat2trans),
    .io_to_pes_6_out_valid(PENetwork_66_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_66_io_to_pes_6_out_bits),
    .io_to_pes_6_sig_stat2trans(PENetwork_66_io_to_pes_6_sig_stat2trans),
    .io_to_pes_7_out_valid(PENetwork_66_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_66_io_to_pes_7_out_bits),
    .io_to_pes_7_sig_stat2trans(PENetwork_66_io_to_pes_7_sig_stat2trans),
    .io_to_pes_8_out_valid(PENetwork_66_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_66_io_to_pes_8_out_bits),
    .io_to_pes_8_sig_stat2trans(PENetwork_66_io_to_pes_8_sig_stat2trans),
    .io_to_pes_9_out_valid(PENetwork_66_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_66_io_to_pes_9_out_bits),
    .io_to_pes_9_sig_stat2trans(PENetwork_66_io_to_pes_9_sig_stat2trans),
    .io_to_pes_10_out_valid(PENetwork_66_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_66_io_to_pes_10_out_bits),
    .io_to_pes_10_sig_stat2trans(PENetwork_66_io_to_pes_10_sig_stat2trans),
    .io_to_pes_11_out_valid(PENetwork_66_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_66_io_to_pes_11_out_bits),
    .io_to_pes_11_sig_stat2trans(PENetwork_66_io_to_pes_11_sig_stat2trans),
    .io_to_pes_12_out_valid(PENetwork_66_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_66_io_to_pes_12_out_bits),
    .io_to_pes_12_sig_stat2trans(PENetwork_66_io_to_pes_12_sig_stat2trans),
    .io_to_pes_13_out_valid(PENetwork_66_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_66_io_to_pes_13_out_bits),
    .io_to_pes_13_sig_stat2trans(PENetwork_66_io_to_pes_13_sig_stat2trans),
    .io_to_pes_14_out_valid(PENetwork_66_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_66_io_to_pes_14_out_bits),
    .io_to_pes_14_sig_stat2trans(PENetwork_66_io_to_pes_14_sig_stat2trans),
    .io_to_pes_15_out_valid(PENetwork_66_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_66_io_to_pes_15_out_bits),
    .io_to_pes_15_sig_stat2trans(PENetwork_66_io_to_pes_15_sig_stat2trans),
    .io_to_pes_16_out_valid(PENetwork_66_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_66_io_to_pes_16_out_bits),
    .io_to_pes_16_sig_stat2trans(PENetwork_66_io_to_pes_16_sig_stat2trans),
    .io_to_pes_17_out_valid(PENetwork_66_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_66_io_to_pes_17_out_bits),
    .io_to_pes_17_sig_stat2trans(PENetwork_66_io_to_pes_17_sig_stat2trans),
    .io_to_pes_18_out_valid(PENetwork_66_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_66_io_to_pes_18_out_bits),
    .io_to_pes_18_sig_stat2trans(PENetwork_66_io_to_pes_18_sig_stat2trans),
    .io_to_pes_19_out_valid(PENetwork_66_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_66_io_to_pes_19_out_bits),
    .io_to_pes_19_sig_stat2trans(PENetwork_66_io_to_pes_19_sig_stat2trans),
    .io_to_pes_20_out_valid(PENetwork_66_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_66_io_to_pes_20_out_bits),
    .io_to_pes_20_sig_stat2trans(PENetwork_66_io_to_pes_20_sig_stat2trans),
    .io_to_pes_21_out_valid(PENetwork_66_io_to_pes_21_out_valid),
    .io_to_pes_21_out_bits(PENetwork_66_io_to_pes_21_out_bits),
    .io_to_pes_21_sig_stat2trans(PENetwork_66_io_to_pes_21_sig_stat2trans),
    .io_to_mem_valid(PENetwork_66_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_66_io_to_mem_bits),
    .io_sig_stat2trans(PENetwork_66_io_sig_stat2trans)
  );
  PENetwork_52 PENetwork_67 ( // @[pe.scala 229:13]
    .clock(PENetwork_67_clock),
    .reset(PENetwork_67_reset),
    .io_to_pes_0_out_valid(PENetwork_67_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_67_io_to_pes_0_out_bits),
    .io_to_pes_0_sig_stat2trans(PENetwork_67_io_to_pes_0_sig_stat2trans),
    .io_to_pes_1_out_valid(PENetwork_67_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_67_io_to_pes_1_out_bits),
    .io_to_pes_1_sig_stat2trans(PENetwork_67_io_to_pes_1_sig_stat2trans),
    .io_to_pes_2_out_valid(PENetwork_67_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_67_io_to_pes_2_out_bits),
    .io_to_pes_2_sig_stat2trans(PENetwork_67_io_to_pes_2_sig_stat2trans),
    .io_to_pes_3_out_valid(PENetwork_67_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_67_io_to_pes_3_out_bits),
    .io_to_pes_3_sig_stat2trans(PENetwork_67_io_to_pes_3_sig_stat2trans),
    .io_to_pes_4_out_valid(PENetwork_67_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_67_io_to_pes_4_out_bits),
    .io_to_pes_4_sig_stat2trans(PENetwork_67_io_to_pes_4_sig_stat2trans),
    .io_to_pes_5_out_valid(PENetwork_67_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_67_io_to_pes_5_out_bits),
    .io_to_pes_5_sig_stat2trans(PENetwork_67_io_to_pes_5_sig_stat2trans),
    .io_to_pes_6_out_valid(PENetwork_67_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_67_io_to_pes_6_out_bits),
    .io_to_pes_6_sig_stat2trans(PENetwork_67_io_to_pes_6_sig_stat2trans),
    .io_to_pes_7_out_valid(PENetwork_67_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_67_io_to_pes_7_out_bits),
    .io_to_pes_7_sig_stat2trans(PENetwork_67_io_to_pes_7_sig_stat2trans),
    .io_to_pes_8_out_valid(PENetwork_67_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_67_io_to_pes_8_out_bits),
    .io_to_pes_8_sig_stat2trans(PENetwork_67_io_to_pes_8_sig_stat2trans),
    .io_to_pes_9_out_valid(PENetwork_67_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_67_io_to_pes_9_out_bits),
    .io_to_pes_9_sig_stat2trans(PENetwork_67_io_to_pes_9_sig_stat2trans),
    .io_to_pes_10_out_valid(PENetwork_67_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_67_io_to_pes_10_out_bits),
    .io_to_pes_10_sig_stat2trans(PENetwork_67_io_to_pes_10_sig_stat2trans),
    .io_to_pes_11_out_valid(PENetwork_67_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_67_io_to_pes_11_out_bits),
    .io_to_pes_11_sig_stat2trans(PENetwork_67_io_to_pes_11_sig_stat2trans),
    .io_to_pes_12_out_valid(PENetwork_67_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_67_io_to_pes_12_out_bits),
    .io_to_pes_12_sig_stat2trans(PENetwork_67_io_to_pes_12_sig_stat2trans),
    .io_to_pes_13_out_valid(PENetwork_67_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_67_io_to_pes_13_out_bits),
    .io_to_pes_13_sig_stat2trans(PENetwork_67_io_to_pes_13_sig_stat2trans),
    .io_to_pes_14_out_valid(PENetwork_67_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_67_io_to_pes_14_out_bits),
    .io_to_pes_14_sig_stat2trans(PENetwork_67_io_to_pes_14_sig_stat2trans),
    .io_to_pes_15_out_valid(PENetwork_67_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_67_io_to_pes_15_out_bits),
    .io_to_pes_15_sig_stat2trans(PENetwork_67_io_to_pes_15_sig_stat2trans),
    .io_to_pes_16_out_valid(PENetwork_67_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_67_io_to_pes_16_out_bits),
    .io_to_pes_16_sig_stat2trans(PENetwork_67_io_to_pes_16_sig_stat2trans),
    .io_to_pes_17_out_valid(PENetwork_67_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_67_io_to_pes_17_out_bits),
    .io_to_pes_17_sig_stat2trans(PENetwork_67_io_to_pes_17_sig_stat2trans),
    .io_to_pes_18_out_valid(PENetwork_67_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_67_io_to_pes_18_out_bits),
    .io_to_pes_18_sig_stat2trans(PENetwork_67_io_to_pes_18_sig_stat2trans),
    .io_to_pes_19_out_valid(PENetwork_67_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_67_io_to_pes_19_out_bits),
    .io_to_pes_19_sig_stat2trans(PENetwork_67_io_to_pes_19_sig_stat2trans),
    .io_to_pes_20_out_valid(PENetwork_67_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_67_io_to_pes_20_out_bits),
    .io_to_pes_20_sig_stat2trans(PENetwork_67_io_to_pes_20_sig_stat2trans),
    .io_to_pes_21_out_valid(PENetwork_67_io_to_pes_21_out_valid),
    .io_to_pes_21_out_bits(PENetwork_67_io_to_pes_21_out_bits),
    .io_to_pes_21_sig_stat2trans(PENetwork_67_io_to_pes_21_sig_stat2trans),
    .io_to_mem_valid(PENetwork_67_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_67_io_to_mem_bits),
    .io_sig_stat2trans(PENetwork_67_io_sig_stat2trans)
  );
  PENetwork_52 PENetwork_68 ( // @[pe.scala 229:13]
    .clock(PENetwork_68_clock),
    .reset(PENetwork_68_reset),
    .io_to_pes_0_out_valid(PENetwork_68_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_68_io_to_pes_0_out_bits),
    .io_to_pes_0_sig_stat2trans(PENetwork_68_io_to_pes_0_sig_stat2trans),
    .io_to_pes_1_out_valid(PENetwork_68_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_68_io_to_pes_1_out_bits),
    .io_to_pes_1_sig_stat2trans(PENetwork_68_io_to_pes_1_sig_stat2trans),
    .io_to_pes_2_out_valid(PENetwork_68_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_68_io_to_pes_2_out_bits),
    .io_to_pes_2_sig_stat2trans(PENetwork_68_io_to_pes_2_sig_stat2trans),
    .io_to_pes_3_out_valid(PENetwork_68_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_68_io_to_pes_3_out_bits),
    .io_to_pes_3_sig_stat2trans(PENetwork_68_io_to_pes_3_sig_stat2trans),
    .io_to_pes_4_out_valid(PENetwork_68_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_68_io_to_pes_4_out_bits),
    .io_to_pes_4_sig_stat2trans(PENetwork_68_io_to_pes_4_sig_stat2trans),
    .io_to_pes_5_out_valid(PENetwork_68_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_68_io_to_pes_5_out_bits),
    .io_to_pes_5_sig_stat2trans(PENetwork_68_io_to_pes_5_sig_stat2trans),
    .io_to_pes_6_out_valid(PENetwork_68_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_68_io_to_pes_6_out_bits),
    .io_to_pes_6_sig_stat2trans(PENetwork_68_io_to_pes_6_sig_stat2trans),
    .io_to_pes_7_out_valid(PENetwork_68_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_68_io_to_pes_7_out_bits),
    .io_to_pes_7_sig_stat2trans(PENetwork_68_io_to_pes_7_sig_stat2trans),
    .io_to_pes_8_out_valid(PENetwork_68_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_68_io_to_pes_8_out_bits),
    .io_to_pes_8_sig_stat2trans(PENetwork_68_io_to_pes_8_sig_stat2trans),
    .io_to_pes_9_out_valid(PENetwork_68_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_68_io_to_pes_9_out_bits),
    .io_to_pes_9_sig_stat2trans(PENetwork_68_io_to_pes_9_sig_stat2trans),
    .io_to_pes_10_out_valid(PENetwork_68_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_68_io_to_pes_10_out_bits),
    .io_to_pes_10_sig_stat2trans(PENetwork_68_io_to_pes_10_sig_stat2trans),
    .io_to_pes_11_out_valid(PENetwork_68_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_68_io_to_pes_11_out_bits),
    .io_to_pes_11_sig_stat2trans(PENetwork_68_io_to_pes_11_sig_stat2trans),
    .io_to_pes_12_out_valid(PENetwork_68_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_68_io_to_pes_12_out_bits),
    .io_to_pes_12_sig_stat2trans(PENetwork_68_io_to_pes_12_sig_stat2trans),
    .io_to_pes_13_out_valid(PENetwork_68_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_68_io_to_pes_13_out_bits),
    .io_to_pes_13_sig_stat2trans(PENetwork_68_io_to_pes_13_sig_stat2trans),
    .io_to_pes_14_out_valid(PENetwork_68_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_68_io_to_pes_14_out_bits),
    .io_to_pes_14_sig_stat2trans(PENetwork_68_io_to_pes_14_sig_stat2trans),
    .io_to_pes_15_out_valid(PENetwork_68_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_68_io_to_pes_15_out_bits),
    .io_to_pes_15_sig_stat2trans(PENetwork_68_io_to_pes_15_sig_stat2trans),
    .io_to_pes_16_out_valid(PENetwork_68_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_68_io_to_pes_16_out_bits),
    .io_to_pes_16_sig_stat2trans(PENetwork_68_io_to_pes_16_sig_stat2trans),
    .io_to_pes_17_out_valid(PENetwork_68_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_68_io_to_pes_17_out_bits),
    .io_to_pes_17_sig_stat2trans(PENetwork_68_io_to_pes_17_sig_stat2trans),
    .io_to_pes_18_out_valid(PENetwork_68_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_68_io_to_pes_18_out_bits),
    .io_to_pes_18_sig_stat2trans(PENetwork_68_io_to_pes_18_sig_stat2trans),
    .io_to_pes_19_out_valid(PENetwork_68_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_68_io_to_pes_19_out_bits),
    .io_to_pes_19_sig_stat2trans(PENetwork_68_io_to_pes_19_sig_stat2trans),
    .io_to_pes_20_out_valid(PENetwork_68_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_68_io_to_pes_20_out_bits),
    .io_to_pes_20_sig_stat2trans(PENetwork_68_io_to_pes_20_sig_stat2trans),
    .io_to_pes_21_out_valid(PENetwork_68_io_to_pes_21_out_valid),
    .io_to_pes_21_out_bits(PENetwork_68_io_to_pes_21_out_bits),
    .io_to_pes_21_sig_stat2trans(PENetwork_68_io_to_pes_21_sig_stat2trans),
    .io_to_mem_valid(PENetwork_68_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_68_io_to_mem_bits),
    .io_sig_stat2trans(PENetwork_68_io_sig_stat2trans)
  );
  PENetwork_52 PENetwork_69 ( // @[pe.scala 229:13]
    .clock(PENetwork_69_clock),
    .reset(PENetwork_69_reset),
    .io_to_pes_0_out_valid(PENetwork_69_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_69_io_to_pes_0_out_bits),
    .io_to_pes_0_sig_stat2trans(PENetwork_69_io_to_pes_0_sig_stat2trans),
    .io_to_pes_1_out_valid(PENetwork_69_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_69_io_to_pes_1_out_bits),
    .io_to_pes_1_sig_stat2trans(PENetwork_69_io_to_pes_1_sig_stat2trans),
    .io_to_pes_2_out_valid(PENetwork_69_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_69_io_to_pes_2_out_bits),
    .io_to_pes_2_sig_stat2trans(PENetwork_69_io_to_pes_2_sig_stat2trans),
    .io_to_pes_3_out_valid(PENetwork_69_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_69_io_to_pes_3_out_bits),
    .io_to_pes_3_sig_stat2trans(PENetwork_69_io_to_pes_3_sig_stat2trans),
    .io_to_pes_4_out_valid(PENetwork_69_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_69_io_to_pes_4_out_bits),
    .io_to_pes_4_sig_stat2trans(PENetwork_69_io_to_pes_4_sig_stat2trans),
    .io_to_pes_5_out_valid(PENetwork_69_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_69_io_to_pes_5_out_bits),
    .io_to_pes_5_sig_stat2trans(PENetwork_69_io_to_pes_5_sig_stat2trans),
    .io_to_pes_6_out_valid(PENetwork_69_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_69_io_to_pes_6_out_bits),
    .io_to_pes_6_sig_stat2trans(PENetwork_69_io_to_pes_6_sig_stat2trans),
    .io_to_pes_7_out_valid(PENetwork_69_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_69_io_to_pes_7_out_bits),
    .io_to_pes_7_sig_stat2trans(PENetwork_69_io_to_pes_7_sig_stat2trans),
    .io_to_pes_8_out_valid(PENetwork_69_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_69_io_to_pes_8_out_bits),
    .io_to_pes_8_sig_stat2trans(PENetwork_69_io_to_pes_8_sig_stat2trans),
    .io_to_pes_9_out_valid(PENetwork_69_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_69_io_to_pes_9_out_bits),
    .io_to_pes_9_sig_stat2trans(PENetwork_69_io_to_pes_9_sig_stat2trans),
    .io_to_pes_10_out_valid(PENetwork_69_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_69_io_to_pes_10_out_bits),
    .io_to_pes_10_sig_stat2trans(PENetwork_69_io_to_pes_10_sig_stat2trans),
    .io_to_pes_11_out_valid(PENetwork_69_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_69_io_to_pes_11_out_bits),
    .io_to_pes_11_sig_stat2trans(PENetwork_69_io_to_pes_11_sig_stat2trans),
    .io_to_pes_12_out_valid(PENetwork_69_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_69_io_to_pes_12_out_bits),
    .io_to_pes_12_sig_stat2trans(PENetwork_69_io_to_pes_12_sig_stat2trans),
    .io_to_pes_13_out_valid(PENetwork_69_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_69_io_to_pes_13_out_bits),
    .io_to_pes_13_sig_stat2trans(PENetwork_69_io_to_pes_13_sig_stat2trans),
    .io_to_pes_14_out_valid(PENetwork_69_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_69_io_to_pes_14_out_bits),
    .io_to_pes_14_sig_stat2trans(PENetwork_69_io_to_pes_14_sig_stat2trans),
    .io_to_pes_15_out_valid(PENetwork_69_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_69_io_to_pes_15_out_bits),
    .io_to_pes_15_sig_stat2trans(PENetwork_69_io_to_pes_15_sig_stat2trans),
    .io_to_pes_16_out_valid(PENetwork_69_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_69_io_to_pes_16_out_bits),
    .io_to_pes_16_sig_stat2trans(PENetwork_69_io_to_pes_16_sig_stat2trans),
    .io_to_pes_17_out_valid(PENetwork_69_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_69_io_to_pes_17_out_bits),
    .io_to_pes_17_sig_stat2trans(PENetwork_69_io_to_pes_17_sig_stat2trans),
    .io_to_pes_18_out_valid(PENetwork_69_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_69_io_to_pes_18_out_bits),
    .io_to_pes_18_sig_stat2trans(PENetwork_69_io_to_pes_18_sig_stat2trans),
    .io_to_pes_19_out_valid(PENetwork_69_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_69_io_to_pes_19_out_bits),
    .io_to_pes_19_sig_stat2trans(PENetwork_69_io_to_pes_19_sig_stat2trans),
    .io_to_pes_20_out_valid(PENetwork_69_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_69_io_to_pes_20_out_bits),
    .io_to_pes_20_sig_stat2trans(PENetwork_69_io_to_pes_20_sig_stat2trans),
    .io_to_pes_21_out_valid(PENetwork_69_io_to_pes_21_out_valid),
    .io_to_pes_21_out_bits(PENetwork_69_io_to_pes_21_out_bits),
    .io_to_pes_21_sig_stat2trans(PENetwork_69_io_to_pes_21_sig_stat2trans),
    .io_to_mem_valid(PENetwork_69_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_69_io_to_mem_bits),
    .io_sig_stat2trans(PENetwork_69_io_sig_stat2trans)
  );
  PENetwork_52 PENetwork_70 ( // @[pe.scala 229:13]
    .clock(PENetwork_70_clock),
    .reset(PENetwork_70_reset),
    .io_to_pes_0_out_valid(PENetwork_70_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_70_io_to_pes_0_out_bits),
    .io_to_pes_0_sig_stat2trans(PENetwork_70_io_to_pes_0_sig_stat2trans),
    .io_to_pes_1_out_valid(PENetwork_70_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_70_io_to_pes_1_out_bits),
    .io_to_pes_1_sig_stat2trans(PENetwork_70_io_to_pes_1_sig_stat2trans),
    .io_to_pes_2_out_valid(PENetwork_70_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_70_io_to_pes_2_out_bits),
    .io_to_pes_2_sig_stat2trans(PENetwork_70_io_to_pes_2_sig_stat2trans),
    .io_to_pes_3_out_valid(PENetwork_70_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_70_io_to_pes_3_out_bits),
    .io_to_pes_3_sig_stat2trans(PENetwork_70_io_to_pes_3_sig_stat2trans),
    .io_to_pes_4_out_valid(PENetwork_70_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_70_io_to_pes_4_out_bits),
    .io_to_pes_4_sig_stat2trans(PENetwork_70_io_to_pes_4_sig_stat2trans),
    .io_to_pes_5_out_valid(PENetwork_70_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_70_io_to_pes_5_out_bits),
    .io_to_pes_5_sig_stat2trans(PENetwork_70_io_to_pes_5_sig_stat2trans),
    .io_to_pes_6_out_valid(PENetwork_70_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_70_io_to_pes_6_out_bits),
    .io_to_pes_6_sig_stat2trans(PENetwork_70_io_to_pes_6_sig_stat2trans),
    .io_to_pes_7_out_valid(PENetwork_70_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_70_io_to_pes_7_out_bits),
    .io_to_pes_7_sig_stat2trans(PENetwork_70_io_to_pes_7_sig_stat2trans),
    .io_to_pes_8_out_valid(PENetwork_70_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_70_io_to_pes_8_out_bits),
    .io_to_pes_8_sig_stat2trans(PENetwork_70_io_to_pes_8_sig_stat2trans),
    .io_to_pes_9_out_valid(PENetwork_70_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_70_io_to_pes_9_out_bits),
    .io_to_pes_9_sig_stat2trans(PENetwork_70_io_to_pes_9_sig_stat2trans),
    .io_to_pes_10_out_valid(PENetwork_70_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_70_io_to_pes_10_out_bits),
    .io_to_pes_10_sig_stat2trans(PENetwork_70_io_to_pes_10_sig_stat2trans),
    .io_to_pes_11_out_valid(PENetwork_70_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_70_io_to_pes_11_out_bits),
    .io_to_pes_11_sig_stat2trans(PENetwork_70_io_to_pes_11_sig_stat2trans),
    .io_to_pes_12_out_valid(PENetwork_70_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_70_io_to_pes_12_out_bits),
    .io_to_pes_12_sig_stat2trans(PENetwork_70_io_to_pes_12_sig_stat2trans),
    .io_to_pes_13_out_valid(PENetwork_70_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_70_io_to_pes_13_out_bits),
    .io_to_pes_13_sig_stat2trans(PENetwork_70_io_to_pes_13_sig_stat2trans),
    .io_to_pes_14_out_valid(PENetwork_70_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_70_io_to_pes_14_out_bits),
    .io_to_pes_14_sig_stat2trans(PENetwork_70_io_to_pes_14_sig_stat2trans),
    .io_to_pes_15_out_valid(PENetwork_70_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_70_io_to_pes_15_out_bits),
    .io_to_pes_15_sig_stat2trans(PENetwork_70_io_to_pes_15_sig_stat2trans),
    .io_to_pes_16_out_valid(PENetwork_70_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_70_io_to_pes_16_out_bits),
    .io_to_pes_16_sig_stat2trans(PENetwork_70_io_to_pes_16_sig_stat2trans),
    .io_to_pes_17_out_valid(PENetwork_70_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_70_io_to_pes_17_out_bits),
    .io_to_pes_17_sig_stat2trans(PENetwork_70_io_to_pes_17_sig_stat2trans),
    .io_to_pes_18_out_valid(PENetwork_70_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_70_io_to_pes_18_out_bits),
    .io_to_pes_18_sig_stat2trans(PENetwork_70_io_to_pes_18_sig_stat2trans),
    .io_to_pes_19_out_valid(PENetwork_70_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_70_io_to_pes_19_out_bits),
    .io_to_pes_19_sig_stat2trans(PENetwork_70_io_to_pes_19_sig_stat2trans),
    .io_to_pes_20_out_valid(PENetwork_70_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_70_io_to_pes_20_out_bits),
    .io_to_pes_20_sig_stat2trans(PENetwork_70_io_to_pes_20_sig_stat2trans),
    .io_to_pes_21_out_valid(PENetwork_70_io_to_pes_21_out_valid),
    .io_to_pes_21_out_bits(PENetwork_70_io_to_pes_21_out_bits),
    .io_to_pes_21_sig_stat2trans(PENetwork_70_io_to_pes_21_sig_stat2trans),
    .io_to_mem_valid(PENetwork_70_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_70_io_to_mem_bits),
    .io_sig_stat2trans(PENetwork_70_io_sig_stat2trans)
  );
  PENetwork_52 PENetwork_71 ( // @[pe.scala 229:13]
    .clock(PENetwork_71_clock),
    .reset(PENetwork_71_reset),
    .io_to_pes_0_out_valid(PENetwork_71_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_71_io_to_pes_0_out_bits),
    .io_to_pes_0_sig_stat2trans(PENetwork_71_io_to_pes_0_sig_stat2trans),
    .io_to_pes_1_out_valid(PENetwork_71_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_71_io_to_pes_1_out_bits),
    .io_to_pes_1_sig_stat2trans(PENetwork_71_io_to_pes_1_sig_stat2trans),
    .io_to_pes_2_out_valid(PENetwork_71_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_71_io_to_pes_2_out_bits),
    .io_to_pes_2_sig_stat2trans(PENetwork_71_io_to_pes_2_sig_stat2trans),
    .io_to_pes_3_out_valid(PENetwork_71_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_71_io_to_pes_3_out_bits),
    .io_to_pes_3_sig_stat2trans(PENetwork_71_io_to_pes_3_sig_stat2trans),
    .io_to_pes_4_out_valid(PENetwork_71_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_71_io_to_pes_4_out_bits),
    .io_to_pes_4_sig_stat2trans(PENetwork_71_io_to_pes_4_sig_stat2trans),
    .io_to_pes_5_out_valid(PENetwork_71_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_71_io_to_pes_5_out_bits),
    .io_to_pes_5_sig_stat2trans(PENetwork_71_io_to_pes_5_sig_stat2trans),
    .io_to_pes_6_out_valid(PENetwork_71_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_71_io_to_pes_6_out_bits),
    .io_to_pes_6_sig_stat2trans(PENetwork_71_io_to_pes_6_sig_stat2trans),
    .io_to_pes_7_out_valid(PENetwork_71_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_71_io_to_pes_7_out_bits),
    .io_to_pes_7_sig_stat2trans(PENetwork_71_io_to_pes_7_sig_stat2trans),
    .io_to_pes_8_out_valid(PENetwork_71_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_71_io_to_pes_8_out_bits),
    .io_to_pes_8_sig_stat2trans(PENetwork_71_io_to_pes_8_sig_stat2trans),
    .io_to_pes_9_out_valid(PENetwork_71_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_71_io_to_pes_9_out_bits),
    .io_to_pes_9_sig_stat2trans(PENetwork_71_io_to_pes_9_sig_stat2trans),
    .io_to_pes_10_out_valid(PENetwork_71_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_71_io_to_pes_10_out_bits),
    .io_to_pes_10_sig_stat2trans(PENetwork_71_io_to_pes_10_sig_stat2trans),
    .io_to_pes_11_out_valid(PENetwork_71_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_71_io_to_pes_11_out_bits),
    .io_to_pes_11_sig_stat2trans(PENetwork_71_io_to_pes_11_sig_stat2trans),
    .io_to_pes_12_out_valid(PENetwork_71_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_71_io_to_pes_12_out_bits),
    .io_to_pes_12_sig_stat2trans(PENetwork_71_io_to_pes_12_sig_stat2trans),
    .io_to_pes_13_out_valid(PENetwork_71_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_71_io_to_pes_13_out_bits),
    .io_to_pes_13_sig_stat2trans(PENetwork_71_io_to_pes_13_sig_stat2trans),
    .io_to_pes_14_out_valid(PENetwork_71_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_71_io_to_pes_14_out_bits),
    .io_to_pes_14_sig_stat2trans(PENetwork_71_io_to_pes_14_sig_stat2trans),
    .io_to_pes_15_out_valid(PENetwork_71_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_71_io_to_pes_15_out_bits),
    .io_to_pes_15_sig_stat2trans(PENetwork_71_io_to_pes_15_sig_stat2trans),
    .io_to_pes_16_out_valid(PENetwork_71_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_71_io_to_pes_16_out_bits),
    .io_to_pes_16_sig_stat2trans(PENetwork_71_io_to_pes_16_sig_stat2trans),
    .io_to_pes_17_out_valid(PENetwork_71_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_71_io_to_pes_17_out_bits),
    .io_to_pes_17_sig_stat2trans(PENetwork_71_io_to_pes_17_sig_stat2trans),
    .io_to_pes_18_out_valid(PENetwork_71_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_71_io_to_pes_18_out_bits),
    .io_to_pes_18_sig_stat2trans(PENetwork_71_io_to_pes_18_sig_stat2trans),
    .io_to_pes_19_out_valid(PENetwork_71_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_71_io_to_pes_19_out_bits),
    .io_to_pes_19_sig_stat2trans(PENetwork_71_io_to_pes_19_sig_stat2trans),
    .io_to_pes_20_out_valid(PENetwork_71_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_71_io_to_pes_20_out_bits),
    .io_to_pes_20_sig_stat2trans(PENetwork_71_io_to_pes_20_sig_stat2trans),
    .io_to_pes_21_out_valid(PENetwork_71_io_to_pes_21_out_valid),
    .io_to_pes_21_out_bits(PENetwork_71_io_to_pes_21_out_bits),
    .io_to_pes_21_sig_stat2trans(PENetwork_71_io_to_pes_21_sig_stat2trans),
    .io_to_mem_valid(PENetwork_71_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_71_io_to_mem_bits),
    .io_sig_stat2trans(PENetwork_71_io_sig_stat2trans)
  );
  PENetwork_52 PENetwork_72 ( // @[pe.scala 229:13]
    .clock(PENetwork_72_clock),
    .reset(PENetwork_72_reset),
    .io_to_pes_0_out_valid(PENetwork_72_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_72_io_to_pes_0_out_bits),
    .io_to_pes_0_sig_stat2trans(PENetwork_72_io_to_pes_0_sig_stat2trans),
    .io_to_pes_1_out_valid(PENetwork_72_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_72_io_to_pes_1_out_bits),
    .io_to_pes_1_sig_stat2trans(PENetwork_72_io_to_pes_1_sig_stat2trans),
    .io_to_pes_2_out_valid(PENetwork_72_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_72_io_to_pes_2_out_bits),
    .io_to_pes_2_sig_stat2trans(PENetwork_72_io_to_pes_2_sig_stat2trans),
    .io_to_pes_3_out_valid(PENetwork_72_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_72_io_to_pes_3_out_bits),
    .io_to_pes_3_sig_stat2trans(PENetwork_72_io_to_pes_3_sig_stat2trans),
    .io_to_pes_4_out_valid(PENetwork_72_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_72_io_to_pes_4_out_bits),
    .io_to_pes_4_sig_stat2trans(PENetwork_72_io_to_pes_4_sig_stat2trans),
    .io_to_pes_5_out_valid(PENetwork_72_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_72_io_to_pes_5_out_bits),
    .io_to_pes_5_sig_stat2trans(PENetwork_72_io_to_pes_5_sig_stat2trans),
    .io_to_pes_6_out_valid(PENetwork_72_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_72_io_to_pes_6_out_bits),
    .io_to_pes_6_sig_stat2trans(PENetwork_72_io_to_pes_6_sig_stat2trans),
    .io_to_pes_7_out_valid(PENetwork_72_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_72_io_to_pes_7_out_bits),
    .io_to_pes_7_sig_stat2trans(PENetwork_72_io_to_pes_7_sig_stat2trans),
    .io_to_pes_8_out_valid(PENetwork_72_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_72_io_to_pes_8_out_bits),
    .io_to_pes_8_sig_stat2trans(PENetwork_72_io_to_pes_8_sig_stat2trans),
    .io_to_pes_9_out_valid(PENetwork_72_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_72_io_to_pes_9_out_bits),
    .io_to_pes_9_sig_stat2trans(PENetwork_72_io_to_pes_9_sig_stat2trans),
    .io_to_pes_10_out_valid(PENetwork_72_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_72_io_to_pes_10_out_bits),
    .io_to_pes_10_sig_stat2trans(PENetwork_72_io_to_pes_10_sig_stat2trans),
    .io_to_pes_11_out_valid(PENetwork_72_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_72_io_to_pes_11_out_bits),
    .io_to_pes_11_sig_stat2trans(PENetwork_72_io_to_pes_11_sig_stat2trans),
    .io_to_pes_12_out_valid(PENetwork_72_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_72_io_to_pes_12_out_bits),
    .io_to_pes_12_sig_stat2trans(PENetwork_72_io_to_pes_12_sig_stat2trans),
    .io_to_pes_13_out_valid(PENetwork_72_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_72_io_to_pes_13_out_bits),
    .io_to_pes_13_sig_stat2trans(PENetwork_72_io_to_pes_13_sig_stat2trans),
    .io_to_pes_14_out_valid(PENetwork_72_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_72_io_to_pes_14_out_bits),
    .io_to_pes_14_sig_stat2trans(PENetwork_72_io_to_pes_14_sig_stat2trans),
    .io_to_pes_15_out_valid(PENetwork_72_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_72_io_to_pes_15_out_bits),
    .io_to_pes_15_sig_stat2trans(PENetwork_72_io_to_pes_15_sig_stat2trans),
    .io_to_pes_16_out_valid(PENetwork_72_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_72_io_to_pes_16_out_bits),
    .io_to_pes_16_sig_stat2trans(PENetwork_72_io_to_pes_16_sig_stat2trans),
    .io_to_pes_17_out_valid(PENetwork_72_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_72_io_to_pes_17_out_bits),
    .io_to_pes_17_sig_stat2trans(PENetwork_72_io_to_pes_17_sig_stat2trans),
    .io_to_pes_18_out_valid(PENetwork_72_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_72_io_to_pes_18_out_bits),
    .io_to_pes_18_sig_stat2trans(PENetwork_72_io_to_pes_18_sig_stat2trans),
    .io_to_pes_19_out_valid(PENetwork_72_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_72_io_to_pes_19_out_bits),
    .io_to_pes_19_sig_stat2trans(PENetwork_72_io_to_pes_19_sig_stat2trans),
    .io_to_pes_20_out_valid(PENetwork_72_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_72_io_to_pes_20_out_bits),
    .io_to_pes_20_sig_stat2trans(PENetwork_72_io_to_pes_20_sig_stat2trans),
    .io_to_pes_21_out_valid(PENetwork_72_io_to_pes_21_out_valid),
    .io_to_pes_21_out_bits(PENetwork_72_io_to_pes_21_out_bits),
    .io_to_pes_21_sig_stat2trans(PENetwork_72_io_to_pes_21_sig_stat2trans),
    .io_to_mem_valid(PENetwork_72_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_72_io_to_mem_bits),
    .io_sig_stat2trans(PENetwork_72_io_sig_stat2trans)
  );
  PENetwork_52 PENetwork_73 ( // @[pe.scala 229:13]
    .clock(PENetwork_73_clock),
    .reset(PENetwork_73_reset),
    .io_to_pes_0_out_valid(PENetwork_73_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_73_io_to_pes_0_out_bits),
    .io_to_pes_0_sig_stat2trans(PENetwork_73_io_to_pes_0_sig_stat2trans),
    .io_to_pes_1_out_valid(PENetwork_73_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_73_io_to_pes_1_out_bits),
    .io_to_pes_1_sig_stat2trans(PENetwork_73_io_to_pes_1_sig_stat2trans),
    .io_to_pes_2_out_valid(PENetwork_73_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_73_io_to_pes_2_out_bits),
    .io_to_pes_2_sig_stat2trans(PENetwork_73_io_to_pes_2_sig_stat2trans),
    .io_to_pes_3_out_valid(PENetwork_73_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_73_io_to_pes_3_out_bits),
    .io_to_pes_3_sig_stat2trans(PENetwork_73_io_to_pes_3_sig_stat2trans),
    .io_to_pes_4_out_valid(PENetwork_73_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_73_io_to_pes_4_out_bits),
    .io_to_pes_4_sig_stat2trans(PENetwork_73_io_to_pes_4_sig_stat2trans),
    .io_to_pes_5_out_valid(PENetwork_73_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_73_io_to_pes_5_out_bits),
    .io_to_pes_5_sig_stat2trans(PENetwork_73_io_to_pes_5_sig_stat2trans),
    .io_to_pes_6_out_valid(PENetwork_73_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_73_io_to_pes_6_out_bits),
    .io_to_pes_6_sig_stat2trans(PENetwork_73_io_to_pes_6_sig_stat2trans),
    .io_to_pes_7_out_valid(PENetwork_73_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_73_io_to_pes_7_out_bits),
    .io_to_pes_7_sig_stat2trans(PENetwork_73_io_to_pes_7_sig_stat2trans),
    .io_to_pes_8_out_valid(PENetwork_73_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_73_io_to_pes_8_out_bits),
    .io_to_pes_8_sig_stat2trans(PENetwork_73_io_to_pes_8_sig_stat2trans),
    .io_to_pes_9_out_valid(PENetwork_73_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_73_io_to_pes_9_out_bits),
    .io_to_pes_9_sig_stat2trans(PENetwork_73_io_to_pes_9_sig_stat2trans),
    .io_to_pes_10_out_valid(PENetwork_73_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_73_io_to_pes_10_out_bits),
    .io_to_pes_10_sig_stat2trans(PENetwork_73_io_to_pes_10_sig_stat2trans),
    .io_to_pes_11_out_valid(PENetwork_73_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_73_io_to_pes_11_out_bits),
    .io_to_pes_11_sig_stat2trans(PENetwork_73_io_to_pes_11_sig_stat2trans),
    .io_to_pes_12_out_valid(PENetwork_73_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_73_io_to_pes_12_out_bits),
    .io_to_pes_12_sig_stat2trans(PENetwork_73_io_to_pes_12_sig_stat2trans),
    .io_to_pes_13_out_valid(PENetwork_73_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_73_io_to_pes_13_out_bits),
    .io_to_pes_13_sig_stat2trans(PENetwork_73_io_to_pes_13_sig_stat2trans),
    .io_to_pes_14_out_valid(PENetwork_73_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_73_io_to_pes_14_out_bits),
    .io_to_pes_14_sig_stat2trans(PENetwork_73_io_to_pes_14_sig_stat2trans),
    .io_to_pes_15_out_valid(PENetwork_73_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_73_io_to_pes_15_out_bits),
    .io_to_pes_15_sig_stat2trans(PENetwork_73_io_to_pes_15_sig_stat2trans),
    .io_to_pes_16_out_valid(PENetwork_73_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_73_io_to_pes_16_out_bits),
    .io_to_pes_16_sig_stat2trans(PENetwork_73_io_to_pes_16_sig_stat2trans),
    .io_to_pes_17_out_valid(PENetwork_73_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_73_io_to_pes_17_out_bits),
    .io_to_pes_17_sig_stat2trans(PENetwork_73_io_to_pes_17_sig_stat2trans),
    .io_to_pes_18_out_valid(PENetwork_73_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_73_io_to_pes_18_out_bits),
    .io_to_pes_18_sig_stat2trans(PENetwork_73_io_to_pes_18_sig_stat2trans),
    .io_to_pes_19_out_valid(PENetwork_73_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_73_io_to_pes_19_out_bits),
    .io_to_pes_19_sig_stat2trans(PENetwork_73_io_to_pes_19_sig_stat2trans),
    .io_to_pes_20_out_valid(PENetwork_73_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_73_io_to_pes_20_out_bits),
    .io_to_pes_20_sig_stat2trans(PENetwork_73_io_to_pes_20_sig_stat2trans),
    .io_to_pes_21_out_valid(PENetwork_73_io_to_pes_21_out_valid),
    .io_to_pes_21_out_bits(PENetwork_73_io_to_pes_21_out_bits),
    .io_to_pes_21_sig_stat2trans(PENetwork_73_io_to_pes_21_sig_stat2trans),
    .io_to_mem_valid(PENetwork_73_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_73_io_to_mem_bits),
    .io_sig_stat2trans(PENetwork_73_io_sig_stat2trans)
  );
  PENetwork_52 PENetwork_74 ( // @[pe.scala 229:13]
    .clock(PENetwork_74_clock),
    .reset(PENetwork_74_reset),
    .io_to_pes_0_out_valid(PENetwork_74_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_74_io_to_pes_0_out_bits),
    .io_to_pes_0_sig_stat2trans(PENetwork_74_io_to_pes_0_sig_stat2trans),
    .io_to_pes_1_out_valid(PENetwork_74_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_74_io_to_pes_1_out_bits),
    .io_to_pes_1_sig_stat2trans(PENetwork_74_io_to_pes_1_sig_stat2trans),
    .io_to_pes_2_out_valid(PENetwork_74_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_74_io_to_pes_2_out_bits),
    .io_to_pes_2_sig_stat2trans(PENetwork_74_io_to_pes_2_sig_stat2trans),
    .io_to_pes_3_out_valid(PENetwork_74_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_74_io_to_pes_3_out_bits),
    .io_to_pes_3_sig_stat2trans(PENetwork_74_io_to_pes_3_sig_stat2trans),
    .io_to_pes_4_out_valid(PENetwork_74_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_74_io_to_pes_4_out_bits),
    .io_to_pes_4_sig_stat2trans(PENetwork_74_io_to_pes_4_sig_stat2trans),
    .io_to_pes_5_out_valid(PENetwork_74_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_74_io_to_pes_5_out_bits),
    .io_to_pes_5_sig_stat2trans(PENetwork_74_io_to_pes_5_sig_stat2trans),
    .io_to_pes_6_out_valid(PENetwork_74_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_74_io_to_pes_6_out_bits),
    .io_to_pes_6_sig_stat2trans(PENetwork_74_io_to_pes_6_sig_stat2trans),
    .io_to_pes_7_out_valid(PENetwork_74_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_74_io_to_pes_7_out_bits),
    .io_to_pes_7_sig_stat2trans(PENetwork_74_io_to_pes_7_sig_stat2trans),
    .io_to_pes_8_out_valid(PENetwork_74_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_74_io_to_pes_8_out_bits),
    .io_to_pes_8_sig_stat2trans(PENetwork_74_io_to_pes_8_sig_stat2trans),
    .io_to_pes_9_out_valid(PENetwork_74_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_74_io_to_pes_9_out_bits),
    .io_to_pes_9_sig_stat2trans(PENetwork_74_io_to_pes_9_sig_stat2trans),
    .io_to_pes_10_out_valid(PENetwork_74_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_74_io_to_pes_10_out_bits),
    .io_to_pes_10_sig_stat2trans(PENetwork_74_io_to_pes_10_sig_stat2trans),
    .io_to_pes_11_out_valid(PENetwork_74_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_74_io_to_pes_11_out_bits),
    .io_to_pes_11_sig_stat2trans(PENetwork_74_io_to_pes_11_sig_stat2trans),
    .io_to_pes_12_out_valid(PENetwork_74_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_74_io_to_pes_12_out_bits),
    .io_to_pes_12_sig_stat2trans(PENetwork_74_io_to_pes_12_sig_stat2trans),
    .io_to_pes_13_out_valid(PENetwork_74_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_74_io_to_pes_13_out_bits),
    .io_to_pes_13_sig_stat2trans(PENetwork_74_io_to_pes_13_sig_stat2trans),
    .io_to_pes_14_out_valid(PENetwork_74_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_74_io_to_pes_14_out_bits),
    .io_to_pes_14_sig_stat2trans(PENetwork_74_io_to_pes_14_sig_stat2trans),
    .io_to_pes_15_out_valid(PENetwork_74_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_74_io_to_pes_15_out_bits),
    .io_to_pes_15_sig_stat2trans(PENetwork_74_io_to_pes_15_sig_stat2trans),
    .io_to_pes_16_out_valid(PENetwork_74_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_74_io_to_pes_16_out_bits),
    .io_to_pes_16_sig_stat2trans(PENetwork_74_io_to_pes_16_sig_stat2trans),
    .io_to_pes_17_out_valid(PENetwork_74_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_74_io_to_pes_17_out_bits),
    .io_to_pes_17_sig_stat2trans(PENetwork_74_io_to_pes_17_sig_stat2trans),
    .io_to_pes_18_out_valid(PENetwork_74_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_74_io_to_pes_18_out_bits),
    .io_to_pes_18_sig_stat2trans(PENetwork_74_io_to_pes_18_sig_stat2trans),
    .io_to_pes_19_out_valid(PENetwork_74_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_74_io_to_pes_19_out_bits),
    .io_to_pes_19_sig_stat2trans(PENetwork_74_io_to_pes_19_sig_stat2trans),
    .io_to_pes_20_out_valid(PENetwork_74_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_74_io_to_pes_20_out_bits),
    .io_to_pes_20_sig_stat2trans(PENetwork_74_io_to_pes_20_sig_stat2trans),
    .io_to_pes_21_out_valid(PENetwork_74_io_to_pes_21_out_valid),
    .io_to_pes_21_out_bits(PENetwork_74_io_to_pes_21_out_bits),
    .io_to_pes_21_sig_stat2trans(PENetwork_74_io_to_pes_21_sig_stat2trans),
    .io_to_mem_valid(PENetwork_74_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_74_io_to_mem_bits),
    .io_sig_stat2trans(PENetwork_74_io_sig_stat2trans)
  );
  PENetwork_52 PENetwork_75 ( // @[pe.scala 229:13]
    .clock(PENetwork_75_clock),
    .reset(PENetwork_75_reset),
    .io_to_pes_0_out_valid(PENetwork_75_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_75_io_to_pes_0_out_bits),
    .io_to_pes_0_sig_stat2trans(PENetwork_75_io_to_pes_0_sig_stat2trans),
    .io_to_pes_1_out_valid(PENetwork_75_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_75_io_to_pes_1_out_bits),
    .io_to_pes_1_sig_stat2trans(PENetwork_75_io_to_pes_1_sig_stat2trans),
    .io_to_pes_2_out_valid(PENetwork_75_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_75_io_to_pes_2_out_bits),
    .io_to_pes_2_sig_stat2trans(PENetwork_75_io_to_pes_2_sig_stat2trans),
    .io_to_pes_3_out_valid(PENetwork_75_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_75_io_to_pes_3_out_bits),
    .io_to_pes_3_sig_stat2trans(PENetwork_75_io_to_pes_3_sig_stat2trans),
    .io_to_pes_4_out_valid(PENetwork_75_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_75_io_to_pes_4_out_bits),
    .io_to_pes_4_sig_stat2trans(PENetwork_75_io_to_pes_4_sig_stat2trans),
    .io_to_pes_5_out_valid(PENetwork_75_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_75_io_to_pes_5_out_bits),
    .io_to_pes_5_sig_stat2trans(PENetwork_75_io_to_pes_5_sig_stat2trans),
    .io_to_pes_6_out_valid(PENetwork_75_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_75_io_to_pes_6_out_bits),
    .io_to_pes_6_sig_stat2trans(PENetwork_75_io_to_pes_6_sig_stat2trans),
    .io_to_pes_7_out_valid(PENetwork_75_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_75_io_to_pes_7_out_bits),
    .io_to_pes_7_sig_stat2trans(PENetwork_75_io_to_pes_7_sig_stat2trans),
    .io_to_pes_8_out_valid(PENetwork_75_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_75_io_to_pes_8_out_bits),
    .io_to_pes_8_sig_stat2trans(PENetwork_75_io_to_pes_8_sig_stat2trans),
    .io_to_pes_9_out_valid(PENetwork_75_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_75_io_to_pes_9_out_bits),
    .io_to_pes_9_sig_stat2trans(PENetwork_75_io_to_pes_9_sig_stat2trans),
    .io_to_pes_10_out_valid(PENetwork_75_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_75_io_to_pes_10_out_bits),
    .io_to_pes_10_sig_stat2trans(PENetwork_75_io_to_pes_10_sig_stat2trans),
    .io_to_pes_11_out_valid(PENetwork_75_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_75_io_to_pes_11_out_bits),
    .io_to_pes_11_sig_stat2trans(PENetwork_75_io_to_pes_11_sig_stat2trans),
    .io_to_pes_12_out_valid(PENetwork_75_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_75_io_to_pes_12_out_bits),
    .io_to_pes_12_sig_stat2trans(PENetwork_75_io_to_pes_12_sig_stat2trans),
    .io_to_pes_13_out_valid(PENetwork_75_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_75_io_to_pes_13_out_bits),
    .io_to_pes_13_sig_stat2trans(PENetwork_75_io_to_pes_13_sig_stat2trans),
    .io_to_pes_14_out_valid(PENetwork_75_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_75_io_to_pes_14_out_bits),
    .io_to_pes_14_sig_stat2trans(PENetwork_75_io_to_pes_14_sig_stat2trans),
    .io_to_pes_15_out_valid(PENetwork_75_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_75_io_to_pes_15_out_bits),
    .io_to_pes_15_sig_stat2trans(PENetwork_75_io_to_pes_15_sig_stat2trans),
    .io_to_pes_16_out_valid(PENetwork_75_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_75_io_to_pes_16_out_bits),
    .io_to_pes_16_sig_stat2trans(PENetwork_75_io_to_pes_16_sig_stat2trans),
    .io_to_pes_17_out_valid(PENetwork_75_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_75_io_to_pes_17_out_bits),
    .io_to_pes_17_sig_stat2trans(PENetwork_75_io_to_pes_17_sig_stat2trans),
    .io_to_pes_18_out_valid(PENetwork_75_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_75_io_to_pes_18_out_bits),
    .io_to_pes_18_sig_stat2trans(PENetwork_75_io_to_pes_18_sig_stat2trans),
    .io_to_pes_19_out_valid(PENetwork_75_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_75_io_to_pes_19_out_bits),
    .io_to_pes_19_sig_stat2trans(PENetwork_75_io_to_pes_19_sig_stat2trans),
    .io_to_pes_20_out_valid(PENetwork_75_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_75_io_to_pes_20_out_bits),
    .io_to_pes_20_sig_stat2trans(PENetwork_75_io_to_pes_20_sig_stat2trans),
    .io_to_pes_21_out_valid(PENetwork_75_io_to_pes_21_out_valid),
    .io_to_pes_21_out_bits(PENetwork_75_io_to_pes_21_out_bits),
    .io_to_pes_21_sig_stat2trans(PENetwork_75_io_to_pes_21_sig_stat2trans),
    .io_to_mem_valid(PENetwork_75_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_75_io_to_mem_bits),
    .io_sig_stat2trans(PENetwork_75_io_sig_stat2trans)
  );
  PENetwork_52 PENetwork_76 ( // @[pe.scala 229:13]
    .clock(PENetwork_76_clock),
    .reset(PENetwork_76_reset),
    .io_to_pes_0_out_valid(PENetwork_76_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_76_io_to_pes_0_out_bits),
    .io_to_pes_0_sig_stat2trans(PENetwork_76_io_to_pes_0_sig_stat2trans),
    .io_to_pes_1_out_valid(PENetwork_76_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_76_io_to_pes_1_out_bits),
    .io_to_pes_1_sig_stat2trans(PENetwork_76_io_to_pes_1_sig_stat2trans),
    .io_to_pes_2_out_valid(PENetwork_76_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_76_io_to_pes_2_out_bits),
    .io_to_pes_2_sig_stat2trans(PENetwork_76_io_to_pes_2_sig_stat2trans),
    .io_to_pes_3_out_valid(PENetwork_76_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_76_io_to_pes_3_out_bits),
    .io_to_pes_3_sig_stat2trans(PENetwork_76_io_to_pes_3_sig_stat2trans),
    .io_to_pes_4_out_valid(PENetwork_76_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_76_io_to_pes_4_out_bits),
    .io_to_pes_4_sig_stat2trans(PENetwork_76_io_to_pes_4_sig_stat2trans),
    .io_to_pes_5_out_valid(PENetwork_76_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_76_io_to_pes_5_out_bits),
    .io_to_pes_5_sig_stat2trans(PENetwork_76_io_to_pes_5_sig_stat2trans),
    .io_to_pes_6_out_valid(PENetwork_76_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_76_io_to_pes_6_out_bits),
    .io_to_pes_6_sig_stat2trans(PENetwork_76_io_to_pes_6_sig_stat2trans),
    .io_to_pes_7_out_valid(PENetwork_76_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_76_io_to_pes_7_out_bits),
    .io_to_pes_7_sig_stat2trans(PENetwork_76_io_to_pes_7_sig_stat2trans),
    .io_to_pes_8_out_valid(PENetwork_76_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_76_io_to_pes_8_out_bits),
    .io_to_pes_8_sig_stat2trans(PENetwork_76_io_to_pes_8_sig_stat2trans),
    .io_to_pes_9_out_valid(PENetwork_76_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_76_io_to_pes_9_out_bits),
    .io_to_pes_9_sig_stat2trans(PENetwork_76_io_to_pes_9_sig_stat2trans),
    .io_to_pes_10_out_valid(PENetwork_76_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_76_io_to_pes_10_out_bits),
    .io_to_pes_10_sig_stat2trans(PENetwork_76_io_to_pes_10_sig_stat2trans),
    .io_to_pes_11_out_valid(PENetwork_76_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_76_io_to_pes_11_out_bits),
    .io_to_pes_11_sig_stat2trans(PENetwork_76_io_to_pes_11_sig_stat2trans),
    .io_to_pes_12_out_valid(PENetwork_76_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_76_io_to_pes_12_out_bits),
    .io_to_pes_12_sig_stat2trans(PENetwork_76_io_to_pes_12_sig_stat2trans),
    .io_to_pes_13_out_valid(PENetwork_76_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_76_io_to_pes_13_out_bits),
    .io_to_pes_13_sig_stat2trans(PENetwork_76_io_to_pes_13_sig_stat2trans),
    .io_to_pes_14_out_valid(PENetwork_76_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_76_io_to_pes_14_out_bits),
    .io_to_pes_14_sig_stat2trans(PENetwork_76_io_to_pes_14_sig_stat2trans),
    .io_to_pes_15_out_valid(PENetwork_76_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_76_io_to_pes_15_out_bits),
    .io_to_pes_15_sig_stat2trans(PENetwork_76_io_to_pes_15_sig_stat2trans),
    .io_to_pes_16_out_valid(PENetwork_76_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_76_io_to_pes_16_out_bits),
    .io_to_pes_16_sig_stat2trans(PENetwork_76_io_to_pes_16_sig_stat2trans),
    .io_to_pes_17_out_valid(PENetwork_76_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_76_io_to_pes_17_out_bits),
    .io_to_pes_17_sig_stat2trans(PENetwork_76_io_to_pes_17_sig_stat2trans),
    .io_to_pes_18_out_valid(PENetwork_76_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_76_io_to_pes_18_out_bits),
    .io_to_pes_18_sig_stat2trans(PENetwork_76_io_to_pes_18_sig_stat2trans),
    .io_to_pes_19_out_valid(PENetwork_76_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_76_io_to_pes_19_out_bits),
    .io_to_pes_19_sig_stat2trans(PENetwork_76_io_to_pes_19_sig_stat2trans),
    .io_to_pes_20_out_valid(PENetwork_76_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_76_io_to_pes_20_out_bits),
    .io_to_pes_20_sig_stat2trans(PENetwork_76_io_to_pes_20_sig_stat2trans),
    .io_to_pes_21_out_valid(PENetwork_76_io_to_pes_21_out_valid),
    .io_to_pes_21_out_bits(PENetwork_76_io_to_pes_21_out_bits),
    .io_to_pes_21_sig_stat2trans(PENetwork_76_io_to_pes_21_sig_stat2trans),
    .io_to_mem_valid(PENetwork_76_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_76_io_to_mem_bits),
    .io_sig_stat2trans(PENetwork_76_io_sig_stat2trans)
  );
  PENetwork_52 PENetwork_77 ( // @[pe.scala 229:13]
    .clock(PENetwork_77_clock),
    .reset(PENetwork_77_reset),
    .io_to_pes_0_out_valid(PENetwork_77_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_77_io_to_pes_0_out_bits),
    .io_to_pes_0_sig_stat2trans(PENetwork_77_io_to_pes_0_sig_stat2trans),
    .io_to_pes_1_out_valid(PENetwork_77_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_77_io_to_pes_1_out_bits),
    .io_to_pes_1_sig_stat2trans(PENetwork_77_io_to_pes_1_sig_stat2trans),
    .io_to_pes_2_out_valid(PENetwork_77_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_77_io_to_pes_2_out_bits),
    .io_to_pes_2_sig_stat2trans(PENetwork_77_io_to_pes_2_sig_stat2trans),
    .io_to_pes_3_out_valid(PENetwork_77_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_77_io_to_pes_3_out_bits),
    .io_to_pes_3_sig_stat2trans(PENetwork_77_io_to_pes_3_sig_stat2trans),
    .io_to_pes_4_out_valid(PENetwork_77_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_77_io_to_pes_4_out_bits),
    .io_to_pes_4_sig_stat2trans(PENetwork_77_io_to_pes_4_sig_stat2trans),
    .io_to_pes_5_out_valid(PENetwork_77_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_77_io_to_pes_5_out_bits),
    .io_to_pes_5_sig_stat2trans(PENetwork_77_io_to_pes_5_sig_stat2trans),
    .io_to_pes_6_out_valid(PENetwork_77_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_77_io_to_pes_6_out_bits),
    .io_to_pes_6_sig_stat2trans(PENetwork_77_io_to_pes_6_sig_stat2trans),
    .io_to_pes_7_out_valid(PENetwork_77_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_77_io_to_pes_7_out_bits),
    .io_to_pes_7_sig_stat2trans(PENetwork_77_io_to_pes_7_sig_stat2trans),
    .io_to_pes_8_out_valid(PENetwork_77_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_77_io_to_pes_8_out_bits),
    .io_to_pes_8_sig_stat2trans(PENetwork_77_io_to_pes_8_sig_stat2trans),
    .io_to_pes_9_out_valid(PENetwork_77_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_77_io_to_pes_9_out_bits),
    .io_to_pes_9_sig_stat2trans(PENetwork_77_io_to_pes_9_sig_stat2trans),
    .io_to_pes_10_out_valid(PENetwork_77_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_77_io_to_pes_10_out_bits),
    .io_to_pes_10_sig_stat2trans(PENetwork_77_io_to_pes_10_sig_stat2trans),
    .io_to_pes_11_out_valid(PENetwork_77_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_77_io_to_pes_11_out_bits),
    .io_to_pes_11_sig_stat2trans(PENetwork_77_io_to_pes_11_sig_stat2trans),
    .io_to_pes_12_out_valid(PENetwork_77_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_77_io_to_pes_12_out_bits),
    .io_to_pes_12_sig_stat2trans(PENetwork_77_io_to_pes_12_sig_stat2trans),
    .io_to_pes_13_out_valid(PENetwork_77_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_77_io_to_pes_13_out_bits),
    .io_to_pes_13_sig_stat2trans(PENetwork_77_io_to_pes_13_sig_stat2trans),
    .io_to_pes_14_out_valid(PENetwork_77_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_77_io_to_pes_14_out_bits),
    .io_to_pes_14_sig_stat2trans(PENetwork_77_io_to_pes_14_sig_stat2trans),
    .io_to_pes_15_out_valid(PENetwork_77_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_77_io_to_pes_15_out_bits),
    .io_to_pes_15_sig_stat2trans(PENetwork_77_io_to_pes_15_sig_stat2trans),
    .io_to_pes_16_out_valid(PENetwork_77_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_77_io_to_pes_16_out_bits),
    .io_to_pes_16_sig_stat2trans(PENetwork_77_io_to_pes_16_sig_stat2trans),
    .io_to_pes_17_out_valid(PENetwork_77_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_77_io_to_pes_17_out_bits),
    .io_to_pes_17_sig_stat2trans(PENetwork_77_io_to_pes_17_sig_stat2trans),
    .io_to_pes_18_out_valid(PENetwork_77_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_77_io_to_pes_18_out_bits),
    .io_to_pes_18_sig_stat2trans(PENetwork_77_io_to_pes_18_sig_stat2trans),
    .io_to_pes_19_out_valid(PENetwork_77_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_77_io_to_pes_19_out_bits),
    .io_to_pes_19_sig_stat2trans(PENetwork_77_io_to_pes_19_sig_stat2trans),
    .io_to_pes_20_out_valid(PENetwork_77_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_77_io_to_pes_20_out_bits),
    .io_to_pes_20_sig_stat2trans(PENetwork_77_io_to_pes_20_sig_stat2trans),
    .io_to_pes_21_out_valid(PENetwork_77_io_to_pes_21_out_valid),
    .io_to_pes_21_out_bits(PENetwork_77_io_to_pes_21_out_bits),
    .io_to_pes_21_sig_stat2trans(PENetwork_77_io_to_pes_21_sig_stat2trans),
    .io_to_mem_valid(PENetwork_77_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_77_io_to_mem_bits),
    .io_sig_stat2trans(PENetwork_77_io_sig_stat2trans)
  );
  PENetwork_52 PENetwork_78 ( // @[pe.scala 229:13]
    .clock(PENetwork_78_clock),
    .reset(PENetwork_78_reset),
    .io_to_pes_0_out_valid(PENetwork_78_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_78_io_to_pes_0_out_bits),
    .io_to_pes_0_sig_stat2trans(PENetwork_78_io_to_pes_0_sig_stat2trans),
    .io_to_pes_1_out_valid(PENetwork_78_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_78_io_to_pes_1_out_bits),
    .io_to_pes_1_sig_stat2trans(PENetwork_78_io_to_pes_1_sig_stat2trans),
    .io_to_pes_2_out_valid(PENetwork_78_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_78_io_to_pes_2_out_bits),
    .io_to_pes_2_sig_stat2trans(PENetwork_78_io_to_pes_2_sig_stat2trans),
    .io_to_pes_3_out_valid(PENetwork_78_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_78_io_to_pes_3_out_bits),
    .io_to_pes_3_sig_stat2trans(PENetwork_78_io_to_pes_3_sig_stat2trans),
    .io_to_pes_4_out_valid(PENetwork_78_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_78_io_to_pes_4_out_bits),
    .io_to_pes_4_sig_stat2trans(PENetwork_78_io_to_pes_4_sig_stat2trans),
    .io_to_pes_5_out_valid(PENetwork_78_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_78_io_to_pes_5_out_bits),
    .io_to_pes_5_sig_stat2trans(PENetwork_78_io_to_pes_5_sig_stat2trans),
    .io_to_pes_6_out_valid(PENetwork_78_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_78_io_to_pes_6_out_bits),
    .io_to_pes_6_sig_stat2trans(PENetwork_78_io_to_pes_6_sig_stat2trans),
    .io_to_pes_7_out_valid(PENetwork_78_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_78_io_to_pes_7_out_bits),
    .io_to_pes_7_sig_stat2trans(PENetwork_78_io_to_pes_7_sig_stat2trans),
    .io_to_pes_8_out_valid(PENetwork_78_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_78_io_to_pes_8_out_bits),
    .io_to_pes_8_sig_stat2trans(PENetwork_78_io_to_pes_8_sig_stat2trans),
    .io_to_pes_9_out_valid(PENetwork_78_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_78_io_to_pes_9_out_bits),
    .io_to_pes_9_sig_stat2trans(PENetwork_78_io_to_pes_9_sig_stat2trans),
    .io_to_pes_10_out_valid(PENetwork_78_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_78_io_to_pes_10_out_bits),
    .io_to_pes_10_sig_stat2trans(PENetwork_78_io_to_pes_10_sig_stat2trans),
    .io_to_pes_11_out_valid(PENetwork_78_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_78_io_to_pes_11_out_bits),
    .io_to_pes_11_sig_stat2trans(PENetwork_78_io_to_pes_11_sig_stat2trans),
    .io_to_pes_12_out_valid(PENetwork_78_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_78_io_to_pes_12_out_bits),
    .io_to_pes_12_sig_stat2trans(PENetwork_78_io_to_pes_12_sig_stat2trans),
    .io_to_pes_13_out_valid(PENetwork_78_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_78_io_to_pes_13_out_bits),
    .io_to_pes_13_sig_stat2trans(PENetwork_78_io_to_pes_13_sig_stat2trans),
    .io_to_pes_14_out_valid(PENetwork_78_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_78_io_to_pes_14_out_bits),
    .io_to_pes_14_sig_stat2trans(PENetwork_78_io_to_pes_14_sig_stat2trans),
    .io_to_pes_15_out_valid(PENetwork_78_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_78_io_to_pes_15_out_bits),
    .io_to_pes_15_sig_stat2trans(PENetwork_78_io_to_pes_15_sig_stat2trans),
    .io_to_pes_16_out_valid(PENetwork_78_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_78_io_to_pes_16_out_bits),
    .io_to_pes_16_sig_stat2trans(PENetwork_78_io_to_pes_16_sig_stat2trans),
    .io_to_pes_17_out_valid(PENetwork_78_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_78_io_to_pes_17_out_bits),
    .io_to_pes_17_sig_stat2trans(PENetwork_78_io_to_pes_17_sig_stat2trans),
    .io_to_pes_18_out_valid(PENetwork_78_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_78_io_to_pes_18_out_bits),
    .io_to_pes_18_sig_stat2trans(PENetwork_78_io_to_pes_18_sig_stat2trans),
    .io_to_pes_19_out_valid(PENetwork_78_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_78_io_to_pes_19_out_bits),
    .io_to_pes_19_sig_stat2trans(PENetwork_78_io_to_pes_19_sig_stat2trans),
    .io_to_pes_20_out_valid(PENetwork_78_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_78_io_to_pes_20_out_bits),
    .io_to_pes_20_sig_stat2trans(PENetwork_78_io_to_pes_20_sig_stat2trans),
    .io_to_pes_21_out_valid(PENetwork_78_io_to_pes_21_out_valid),
    .io_to_pes_21_out_bits(PENetwork_78_io_to_pes_21_out_bits),
    .io_to_pes_21_sig_stat2trans(PENetwork_78_io_to_pes_21_sig_stat2trans),
    .io_to_mem_valid(PENetwork_78_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_78_io_to_mem_bits),
    .io_sig_stat2trans(PENetwork_78_io_sig_stat2trans)
  );
  PENetwork_52 PENetwork_79 ( // @[pe.scala 229:13]
    .clock(PENetwork_79_clock),
    .reset(PENetwork_79_reset),
    .io_to_pes_0_out_valid(PENetwork_79_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_79_io_to_pes_0_out_bits),
    .io_to_pes_0_sig_stat2trans(PENetwork_79_io_to_pes_0_sig_stat2trans),
    .io_to_pes_1_out_valid(PENetwork_79_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_79_io_to_pes_1_out_bits),
    .io_to_pes_1_sig_stat2trans(PENetwork_79_io_to_pes_1_sig_stat2trans),
    .io_to_pes_2_out_valid(PENetwork_79_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_79_io_to_pes_2_out_bits),
    .io_to_pes_2_sig_stat2trans(PENetwork_79_io_to_pes_2_sig_stat2trans),
    .io_to_pes_3_out_valid(PENetwork_79_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_79_io_to_pes_3_out_bits),
    .io_to_pes_3_sig_stat2trans(PENetwork_79_io_to_pes_3_sig_stat2trans),
    .io_to_pes_4_out_valid(PENetwork_79_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_79_io_to_pes_4_out_bits),
    .io_to_pes_4_sig_stat2trans(PENetwork_79_io_to_pes_4_sig_stat2trans),
    .io_to_pes_5_out_valid(PENetwork_79_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_79_io_to_pes_5_out_bits),
    .io_to_pes_5_sig_stat2trans(PENetwork_79_io_to_pes_5_sig_stat2trans),
    .io_to_pes_6_out_valid(PENetwork_79_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_79_io_to_pes_6_out_bits),
    .io_to_pes_6_sig_stat2trans(PENetwork_79_io_to_pes_6_sig_stat2trans),
    .io_to_pes_7_out_valid(PENetwork_79_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_79_io_to_pes_7_out_bits),
    .io_to_pes_7_sig_stat2trans(PENetwork_79_io_to_pes_7_sig_stat2trans),
    .io_to_pes_8_out_valid(PENetwork_79_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_79_io_to_pes_8_out_bits),
    .io_to_pes_8_sig_stat2trans(PENetwork_79_io_to_pes_8_sig_stat2trans),
    .io_to_pes_9_out_valid(PENetwork_79_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_79_io_to_pes_9_out_bits),
    .io_to_pes_9_sig_stat2trans(PENetwork_79_io_to_pes_9_sig_stat2trans),
    .io_to_pes_10_out_valid(PENetwork_79_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_79_io_to_pes_10_out_bits),
    .io_to_pes_10_sig_stat2trans(PENetwork_79_io_to_pes_10_sig_stat2trans),
    .io_to_pes_11_out_valid(PENetwork_79_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_79_io_to_pes_11_out_bits),
    .io_to_pes_11_sig_stat2trans(PENetwork_79_io_to_pes_11_sig_stat2trans),
    .io_to_pes_12_out_valid(PENetwork_79_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_79_io_to_pes_12_out_bits),
    .io_to_pes_12_sig_stat2trans(PENetwork_79_io_to_pes_12_sig_stat2trans),
    .io_to_pes_13_out_valid(PENetwork_79_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_79_io_to_pes_13_out_bits),
    .io_to_pes_13_sig_stat2trans(PENetwork_79_io_to_pes_13_sig_stat2trans),
    .io_to_pes_14_out_valid(PENetwork_79_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_79_io_to_pes_14_out_bits),
    .io_to_pes_14_sig_stat2trans(PENetwork_79_io_to_pes_14_sig_stat2trans),
    .io_to_pes_15_out_valid(PENetwork_79_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_79_io_to_pes_15_out_bits),
    .io_to_pes_15_sig_stat2trans(PENetwork_79_io_to_pes_15_sig_stat2trans),
    .io_to_pes_16_out_valid(PENetwork_79_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_79_io_to_pes_16_out_bits),
    .io_to_pes_16_sig_stat2trans(PENetwork_79_io_to_pes_16_sig_stat2trans),
    .io_to_pes_17_out_valid(PENetwork_79_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_79_io_to_pes_17_out_bits),
    .io_to_pes_17_sig_stat2trans(PENetwork_79_io_to_pes_17_sig_stat2trans),
    .io_to_pes_18_out_valid(PENetwork_79_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_79_io_to_pes_18_out_bits),
    .io_to_pes_18_sig_stat2trans(PENetwork_79_io_to_pes_18_sig_stat2trans),
    .io_to_pes_19_out_valid(PENetwork_79_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_79_io_to_pes_19_out_bits),
    .io_to_pes_19_sig_stat2trans(PENetwork_79_io_to_pes_19_sig_stat2trans),
    .io_to_pes_20_out_valid(PENetwork_79_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_79_io_to_pes_20_out_bits),
    .io_to_pes_20_sig_stat2trans(PENetwork_79_io_to_pes_20_sig_stat2trans),
    .io_to_pes_21_out_valid(PENetwork_79_io_to_pes_21_out_valid),
    .io_to_pes_21_out_bits(PENetwork_79_io_to_pes_21_out_bits),
    .io_to_pes_21_sig_stat2trans(PENetwork_79_io_to_pes_21_sig_stat2trans),
    .io_to_mem_valid(PENetwork_79_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_79_io_to_mem_bits),
    .io_sig_stat2trans(PENetwork_79_io_sig_stat2trans)
  );
  PENetwork_52 PENetwork_80 ( // @[pe.scala 229:13]
    .clock(PENetwork_80_clock),
    .reset(PENetwork_80_reset),
    .io_to_pes_0_out_valid(PENetwork_80_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_80_io_to_pes_0_out_bits),
    .io_to_pes_0_sig_stat2trans(PENetwork_80_io_to_pes_0_sig_stat2trans),
    .io_to_pes_1_out_valid(PENetwork_80_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_80_io_to_pes_1_out_bits),
    .io_to_pes_1_sig_stat2trans(PENetwork_80_io_to_pes_1_sig_stat2trans),
    .io_to_pes_2_out_valid(PENetwork_80_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_80_io_to_pes_2_out_bits),
    .io_to_pes_2_sig_stat2trans(PENetwork_80_io_to_pes_2_sig_stat2trans),
    .io_to_pes_3_out_valid(PENetwork_80_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_80_io_to_pes_3_out_bits),
    .io_to_pes_3_sig_stat2trans(PENetwork_80_io_to_pes_3_sig_stat2trans),
    .io_to_pes_4_out_valid(PENetwork_80_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_80_io_to_pes_4_out_bits),
    .io_to_pes_4_sig_stat2trans(PENetwork_80_io_to_pes_4_sig_stat2trans),
    .io_to_pes_5_out_valid(PENetwork_80_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_80_io_to_pes_5_out_bits),
    .io_to_pes_5_sig_stat2trans(PENetwork_80_io_to_pes_5_sig_stat2trans),
    .io_to_pes_6_out_valid(PENetwork_80_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_80_io_to_pes_6_out_bits),
    .io_to_pes_6_sig_stat2trans(PENetwork_80_io_to_pes_6_sig_stat2trans),
    .io_to_pes_7_out_valid(PENetwork_80_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_80_io_to_pes_7_out_bits),
    .io_to_pes_7_sig_stat2trans(PENetwork_80_io_to_pes_7_sig_stat2trans),
    .io_to_pes_8_out_valid(PENetwork_80_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_80_io_to_pes_8_out_bits),
    .io_to_pes_8_sig_stat2trans(PENetwork_80_io_to_pes_8_sig_stat2trans),
    .io_to_pes_9_out_valid(PENetwork_80_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_80_io_to_pes_9_out_bits),
    .io_to_pes_9_sig_stat2trans(PENetwork_80_io_to_pes_9_sig_stat2trans),
    .io_to_pes_10_out_valid(PENetwork_80_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_80_io_to_pes_10_out_bits),
    .io_to_pes_10_sig_stat2trans(PENetwork_80_io_to_pes_10_sig_stat2trans),
    .io_to_pes_11_out_valid(PENetwork_80_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_80_io_to_pes_11_out_bits),
    .io_to_pes_11_sig_stat2trans(PENetwork_80_io_to_pes_11_sig_stat2trans),
    .io_to_pes_12_out_valid(PENetwork_80_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_80_io_to_pes_12_out_bits),
    .io_to_pes_12_sig_stat2trans(PENetwork_80_io_to_pes_12_sig_stat2trans),
    .io_to_pes_13_out_valid(PENetwork_80_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_80_io_to_pes_13_out_bits),
    .io_to_pes_13_sig_stat2trans(PENetwork_80_io_to_pes_13_sig_stat2trans),
    .io_to_pes_14_out_valid(PENetwork_80_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_80_io_to_pes_14_out_bits),
    .io_to_pes_14_sig_stat2trans(PENetwork_80_io_to_pes_14_sig_stat2trans),
    .io_to_pes_15_out_valid(PENetwork_80_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_80_io_to_pes_15_out_bits),
    .io_to_pes_15_sig_stat2trans(PENetwork_80_io_to_pes_15_sig_stat2trans),
    .io_to_pes_16_out_valid(PENetwork_80_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_80_io_to_pes_16_out_bits),
    .io_to_pes_16_sig_stat2trans(PENetwork_80_io_to_pes_16_sig_stat2trans),
    .io_to_pes_17_out_valid(PENetwork_80_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_80_io_to_pes_17_out_bits),
    .io_to_pes_17_sig_stat2trans(PENetwork_80_io_to_pes_17_sig_stat2trans),
    .io_to_pes_18_out_valid(PENetwork_80_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_80_io_to_pes_18_out_bits),
    .io_to_pes_18_sig_stat2trans(PENetwork_80_io_to_pes_18_sig_stat2trans),
    .io_to_pes_19_out_valid(PENetwork_80_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_80_io_to_pes_19_out_bits),
    .io_to_pes_19_sig_stat2trans(PENetwork_80_io_to_pes_19_sig_stat2trans),
    .io_to_pes_20_out_valid(PENetwork_80_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_80_io_to_pes_20_out_bits),
    .io_to_pes_20_sig_stat2trans(PENetwork_80_io_to_pes_20_sig_stat2trans),
    .io_to_pes_21_out_valid(PENetwork_80_io_to_pes_21_out_valid),
    .io_to_pes_21_out_bits(PENetwork_80_io_to_pes_21_out_bits),
    .io_to_pes_21_sig_stat2trans(PENetwork_80_io_to_pes_21_sig_stat2trans),
    .io_to_mem_valid(PENetwork_80_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_80_io_to_mem_bits),
    .io_sig_stat2trans(PENetwork_80_io_sig_stat2trans)
  );
  PENetwork_52 PENetwork_81 ( // @[pe.scala 229:13]
    .clock(PENetwork_81_clock),
    .reset(PENetwork_81_reset),
    .io_to_pes_0_out_valid(PENetwork_81_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_81_io_to_pes_0_out_bits),
    .io_to_pes_0_sig_stat2trans(PENetwork_81_io_to_pes_0_sig_stat2trans),
    .io_to_pes_1_out_valid(PENetwork_81_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_81_io_to_pes_1_out_bits),
    .io_to_pes_1_sig_stat2trans(PENetwork_81_io_to_pes_1_sig_stat2trans),
    .io_to_pes_2_out_valid(PENetwork_81_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_81_io_to_pes_2_out_bits),
    .io_to_pes_2_sig_stat2trans(PENetwork_81_io_to_pes_2_sig_stat2trans),
    .io_to_pes_3_out_valid(PENetwork_81_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_81_io_to_pes_3_out_bits),
    .io_to_pes_3_sig_stat2trans(PENetwork_81_io_to_pes_3_sig_stat2trans),
    .io_to_pes_4_out_valid(PENetwork_81_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_81_io_to_pes_4_out_bits),
    .io_to_pes_4_sig_stat2trans(PENetwork_81_io_to_pes_4_sig_stat2trans),
    .io_to_pes_5_out_valid(PENetwork_81_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_81_io_to_pes_5_out_bits),
    .io_to_pes_5_sig_stat2trans(PENetwork_81_io_to_pes_5_sig_stat2trans),
    .io_to_pes_6_out_valid(PENetwork_81_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_81_io_to_pes_6_out_bits),
    .io_to_pes_6_sig_stat2trans(PENetwork_81_io_to_pes_6_sig_stat2trans),
    .io_to_pes_7_out_valid(PENetwork_81_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_81_io_to_pes_7_out_bits),
    .io_to_pes_7_sig_stat2trans(PENetwork_81_io_to_pes_7_sig_stat2trans),
    .io_to_pes_8_out_valid(PENetwork_81_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_81_io_to_pes_8_out_bits),
    .io_to_pes_8_sig_stat2trans(PENetwork_81_io_to_pes_8_sig_stat2trans),
    .io_to_pes_9_out_valid(PENetwork_81_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_81_io_to_pes_9_out_bits),
    .io_to_pes_9_sig_stat2trans(PENetwork_81_io_to_pes_9_sig_stat2trans),
    .io_to_pes_10_out_valid(PENetwork_81_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_81_io_to_pes_10_out_bits),
    .io_to_pes_10_sig_stat2trans(PENetwork_81_io_to_pes_10_sig_stat2trans),
    .io_to_pes_11_out_valid(PENetwork_81_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_81_io_to_pes_11_out_bits),
    .io_to_pes_11_sig_stat2trans(PENetwork_81_io_to_pes_11_sig_stat2trans),
    .io_to_pes_12_out_valid(PENetwork_81_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_81_io_to_pes_12_out_bits),
    .io_to_pes_12_sig_stat2trans(PENetwork_81_io_to_pes_12_sig_stat2trans),
    .io_to_pes_13_out_valid(PENetwork_81_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_81_io_to_pes_13_out_bits),
    .io_to_pes_13_sig_stat2trans(PENetwork_81_io_to_pes_13_sig_stat2trans),
    .io_to_pes_14_out_valid(PENetwork_81_io_to_pes_14_out_valid),
    .io_to_pes_14_out_bits(PENetwork_81_io_to_pes_14_out_bits),
    .io_to_pes_14_sig_stat2trans(PENetwork_81_io_to_pes_14_sig_stat2trans),
    .io_to_pes_15_out_valid(PENetwork_81_io_to_pes_15_out_valid),
    .io_to_pes_15_out_bits(PENetwork_81_io_to_pes_15_out_bits),
    .io_to_pes_15_sig_stat2trans(PENetwork_81_io_to_pes_15_sig_stat2trans),
    .io_to_pes_16_out_valid(PENetwork_81_io_to_pes_16_out_valid),
    .io_to_pes_16_out_bits(PENetwork_81_io_to_pes_16_out_bits),
    .io_to_pes_16_sig_stat2trans(PENetwork_81_io_to_pes_16_sig_stat2trans),
    .io_to_pes_17_out_valid(PENetwork_81_io_to_pes_17_out_valid),
    .io_to_pes_17_out_bits(PENetwork_81_io_to_pes_17_out_bits),
    .io_to_pes_17_sig_stat2trans(PENetwork_81_io_to_pes_17_sig_stat2trans),
    .io_to_pes_18_out_valid(PENetwork_81_io_to_pes_18_out_valid),
    .io_to_pes_18_out_bits(PENetwork_81_io_to_pes_18_out_bits),
    .io_to_pes_18_sig_stat2trans(PENetwork_81_io_to_pes_18_sig_stat2trans),
    .io_to_pes_19_out_valid(PENetwork_81_io_to_pes_19_out_valid),
    .io_to_pes_19_out_bits(PENetwork_81_io_to_pes_19_out_bits),
    .io_to_pes_19_sig_stat2trans(PENetwork_81_io_to_pes_19_sig_stat2trans),
    .io_to_pes_20_out_valid(PENetwork_81_io_to_pes_20_out_valid),
    .io_to_pes_20_out_bits(PENetwork_81_io_to_pes_20_out_bits),
    .io_to_pes_20_sig_stat2trans(PENetwork_81_io_to_pes_20_sig_stat2trans),
    .io_to_pes_21_out_valid(PENetwork_81_io_to_pes_21_out_valid),
    .io_to_pes_21_out_bits(PENetwork_81_io_to_pes_21_out_bits),
    .io_to_pes_21_sig_stat2trans(PENetwork_81_io_to_pes_21_sig_stat2trans),
    .io_to_mem_valid(PENetwork_81_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_81_io_to_mem_bits),
    .io_sig_stat2trans(PENetwork_81_io_sig_stat2trans)
  );
  MemController MemController ( // @[pe.scala 303:15]
    .clock(MemController_clock),
    .reset(MemController_reset),
    .io_rd_valid(MemController_io_rd_valid),
    .io_wr_valid(MemController_io_wr_valid),
    .io_rd_data_valid(MemController_io_rd_data_valid),
    .io_rd_data_bits(MemController_io_rd_data_bits),
    .io_wr_data_valid(MemController_io_wr_data_valid),
    .io_wr_data_bits(MemController_io_wr_data_bits)
  );
  MemController MemController_1 ( // @[pe.scala 303:15]
    .clock(MemController_1_clock),
    .reset(MemController_1_reset),
    .io_rd_valid(MemController_1_io_rd_valid),
    .io_wr_valid(MemController_1_io_wr_valid),
    .io_rd_data_valid(MemController_1_io_rd_data_valid),
    .io_rd_data_bits(MemController_1_io_rd_data_bits),
    .io_wr_data_valid(MemController_1_io_wr_data_valid),
    .io_wr_data_bits(MemController_1_io_wr_data_bits)
  );
  MemController MemController_2 ( // @[pe.scala 303:15]
    .clock(MemController_2_clock),
    .reset(MemController_2_reset),
    .io_rd_valid(MemController_2_io_rd_valid),
    .io_wr_valid(MemController_2_io_wr_valid),
    .io_rd_data_valid(MemController_2_io_rd_data_valid),
    .io_rd_data_bits(MemController_2_io_rd_data_bits),
    .io_wr_data_valid(MemController_2_io_wr_data_valid),
    .io_wr_data_bits(MemController_2_io_wr_data_bits)
  );
  MemController MemController_3 ( // @[pe.scala 303:15]
    .clock(MemController_3_clock),
    .reset(MemController_3_reset),
    .io_rd_valid(MemController_3_io_rd_valid),
    .io_wr_valid(MemController_3_io_wr_valid),
    .io_rd_data_valid(MemController_3_io_rd_data_valid),
    .io_rd_data_bits(MemController_3_io_rd_data_bits),
    .io_wr_data_valid(MemController_3_io_wr_data_valid),
    .io_wr_data_bits(MemController_3_io_wr_data_bits)
  );
  MemController MemController_4 ( // @[pe.scala 303:15]
    .clock(MemController_4_clock),
    .reset(MemController_4_reset),
    .io_rd_valid(MemController_4_io_rd_valid),
    .io_wr_valid(MemController_4_io_wr_valid),
    .io_rd_data_valid(MemController_4_io_rd_data_valid),
    .io_rd_data_bits(MemController_4_io_rd_data_bits),
    .io_wr_data_valid(MemController_4_io_wr_data_valid),
    .io_wr_data_bits(MemController_4_io_wr_data_bits)
  );
  MemController MemController_5 ( // @[pe.scala 303:15]
    .clock(MemController_5_clock),
    .reset(MemController_5_reset),
    .io_rd_valid(MemController_5_io_rd_valid),
    .io_wr_valid(MemController_5_io_wr_valid),
    .io_rd_data_valid(MemController_5_io_rd_data_valid),
    .io_rd_data_bits(MemController_5_io_rd_data_bits),
    .io_wr_data_valid(MemController_5_io_wr_data_valid),
    .io_wr_data_bits(MemController_5_io_wr_data_bits)
  );
  MemController MemController_6 ( // @[pe.scala 303:15]
    .clock(MemController_6_clock),
    .reset(MemController_6_reset),
    .io_rd_valid(MemController_6_io_rd_valid),
    .io_wr_valid(MemController_6_io_wr_valid),
    .io_rd_data_valid(MemController_6_io_rd_data_valid),
    .io_rd_data_bits(MemController_6_io_rd_data_bits),
    .io_wr_data_valid(MemController_6_io_wr_data_valid),
    .io_wr_data_bits(MemController_6_io_wr_data_bits)
  );
  MemController MemController_7 ( // @[pe.scala 303:15]
    .clock(MemController_7_clock),
    .reset(MemController_7_reset),
    .io_rd_valid(MemController_7_io_rd_valid),
    .io_wr_valid(MemController_7_io_wr_valid),
    .io_rd_data_valid(MemController_7_io_rd_data_valid),
    .io_rd_data_bits(MemController_7_io_rd_data_bits),
    .io_wr_data_valid(MemController_7_io_wr_data_valid),
    .io_wr_data_bits(MemController_7_io_wr_data_bits)
  );
  MemController MemController_8 ( // @[pe.scala 303:15]
    .clock(MemController_8_clock),
    .reset(MemController_8_reset),
    .io_rd_valid(MemController_8_io_rd_valid),
    .io_wr_valid(MemController_8_io_wr_valid),
    .io_rd_data_valid(MemController_8_io_rd_data_valid),
    .io_rd_data_bits(MemController_8_io_rd_data_bits),
    .io_wr_data_valid(MemController_8_io_wr_data_valid),
    .io_wr_data_bits(MemController_8_io_wr_data_bits)
  );
  MemController MemController_9 ( // @[pe.scala 303:15]
    .clock(MemController_9_clock),
    .reset(MemController_9_reset),
    .io_rd_valid(MemController_9_io_rd_valid),
    .io_wr_valid(MemController_9_io_wr_valid),
    .io_rd_data_valid(MemController_9_io_rd_data_valid),
    .io_rd_data_bits(MemController_9_io_rd_data_bits),
    .io_wr_data_valid(MemController_9_io_wr_data_valid),
    .io_wr_data_bits(MemController_9_io_wr_data_bits)
  );
  MemController MemController_10 ( // @[pe.scala 303:15]
    .clock(MemController_10_clock),
    .reset(MemController_10_reset),
    .io_rd_valid(MemController_10_io_rd_valid),
    .io_wr_valid(MemController_10_io_wr_valid),
    .io_rd_data_valid(MemController_10_io_rd_data_valid),
    .io_rd_data_bits(MemController_10_io_rd_data_bits),
    .io_wr_data_valid(MemController_10_io_wr_data_valid),
    .io_wr_data_bits(MemController_10_io_wr_data_bits)
  );
  MemController MemController_11 ( // @[pe.scala 303:15]
    .clock(MemController_11_clock),
    .reset(MemController_11_reset),
    .io_rd_valid(MemController_11_io_rd_valid),
    .io_wr_valid(MemController_11_io_wr_valid),
    .io_rd_data_valid(MemController_11_io_rd_data_valid),
    .io_rd_data_bits(MemController_11_io_rd_data_bits),
    .io_wr_data_valid(MemController_11_io_wr_data_valid),
    .io_wr_data_bits(MemController_11_io_wr_data_bits)
  );
  MemController MemController_12 ( // @[pe.scala 303:15]
    .clock(MemController_12_clock),
    .reset(MemController_12_reset),
    .io_rd_valid(MemController_12_io_rd_valid),
    .io_wr_valid(MemController_12_io_wr_valid),
    .io_rd_data_valid(MemController_12_io_rd_data_valid),
    .io_rd_data_bits(MemController_12_io_rd_data_bits),
    .io_wr_data_valid(MemController_12_io_wr_data_valid),
    .io_wr_data_bits(MemController_12_io_wr_data_bits)
  );
  MemController MemController_13 ( // @[pe.scala 303:15]
    .clock(MemController_13_clock),
    .reset(MemController_13_reset),
    .io_rd_valid(MemController_13_io_rd_valid),
    .io_wr_valid(MemController_13_io_wr_valid),
    .io_rd_data_valid(MemController_13_io_rd_data_valid),
    .io_rd_data_bits(MemController_13_io_rd_data_bits),
    .io_wr_data_valid(MemController_13_io_wr_data_valid),
    .io_wr_data_bits(MemController_13_io_wr_data_bits)
  );
  MemController MemController_14 ( // @[pe.scala 303:15]
    .clock(MemController_14_clock),
    .reset(MemController_14_reset),
    .io_rd_valid(MemController_14_io_rd_valid),
    .io_wr_valid(MemController_14_io_wr_valid),
    .io_rd_data_valid(MemController_14_io_rd_data_valid),
    .io_rd_data_bits(MemController_14_io_rd_data_bits),
    .io_wr_data_valid(MemController_14_io_wr_data_valid),
    .io_wr_data_bits(MemController_14_io_wr_data_bits)
  );
  MemController MemController_15 ( // @[pe.scala 303:15]
    .clock(MemController_15_clock),
    .reset(MemController_15_reset),
    .io_rd_valid(MemController_15_io_rd_valid),
    .io_wr_valid(MemController_15_io_wr_valid),
    .io_rd_data_valid(MemController_15_io_rd_data_valid),
    .io_rd_data_bits(MemController_15_io_rd_data_bits),
    .io_wr_data_valid(MemController_15_io_wr_data_valid),
    .io_wr_data_bits(MemController_15_io_wr_data_bits)
  );
  MemController MemController_16 ( // @[pe.scala 303:15]
    .clock(MemController_16_clock),
    .reset(MemController_16_reset),
    .io_rd_valid(MemController_16_io_rd_valid),
    .io_wr_valid(MemController_16_io_wr_valid),
    .io_rd_data_valid(MemController_16_io_rd_data_valid),
    .io_rd_data_bits(MemController_16_io_rd_data_bits),
    .io_wr_data_valid(MemController_16_io_wr_data_valid),
    .io_wr_data_bits(MemController_16_io_wr_data_bits)
  );
  MemController MemController_17 ( // @[pe.scala 303:15]
    .clock(MemController_17_clock),
    .reset(MemController_17_reset),
    .io_rd_valid(MemController_17_io_rd_valid),
    .io_wr_valid(MemController_17_io_wr_valid),
    .io_rd_data_valid(MemController_17_io_rd_data_valid),
    .io_rd_data_bits(MemController_17_io_rd_data_bits),
    .io_wr_data_valid(MemController_17_io_wr_data_valid),
    .io_wr_data_bits(MemController_17_io_wr_data_bits)
  );
  MemController MemController_18 ( // @[pe.scala 303:15]
    .clock(MemController_18_clock),
    .reset(MemController_18_reset),
    .io_rd_valid(MemController_18_io_rd_valid),
    .io_wr_valid(MemController_18_io_wr_valid),
    .io_rd_data_valid(MemController_18_io_rd_data_valid),
    .io_rd_data_bits(MemController_18_io_rd_data_bits),
    .io_wr_data_valid(MemController_18_io_wr_data_valid),
    .io_wr_data_bits(MemController_18_io_wr_data_bits)
  );
  MemController MemController_19 ( // @[pe.scala 303:15]
    .clock(MemController_19_clock),
    .reset(MemController_19_reset),
    .io_rd_valid(MemController_19_io_rd_valid),
    .io_wr_valid(MemController_19_io_wr_valid),
    .io_rd_data_valid(MemController_19_io_rd_data_valid),
    .io_rd_data_bits(MemController_19_io_rd_data_bits),
    .io_wr_data_valid(MemController_19_io_wr_data_valid),
    .io_wr_data_bits(MemController_19_io_wr_data_bits)
  );
  MemController MemController_20 ( // @[pe.scala 303:15]
    .clock(MemController_20_clock),
    .reset(MemController_20_reset),
    .io_rd_valid(MemController_20_io_rd_valid),
    .io_wr_valid(MemController_20_io_wr_valid),
    .io_rd_data_valid(MemController_20_io_rd_data_valid),
    .io_rd_data_bits(MemController_20_io_rd_data_bits),
    .io_wr_data_valid(MemController_20_io_wr_data_valid),
    .io_wr_data_bits(MemController_20_io_wr_data_bits)
  );
  MemController MemController_21 ( // @[pe.scala 303:15]
    .clock(MemController_21_clock),
    .reset(MemController_21_reset),
    .io_rd_valid(MemController_21_io_rd_valid),
    .io_wr_valid(MemController_21_io_wr_valid),
    .io_rd_data_valid(MemController_21_io_rd_data_valid),
    .io_rd_data_bits(MemController_21_io_rd_data_bits),
    .io_wr_data_valid(MemController_21_io_wr_data_valid),
    .io_wr_data_bits(MemController_21_io_wr_data_bits)
  );
  MemController_22 MemController_22 ( // @[pe.scala 303:15]
    .clock(MemController_22_clock),
    .reset(MemController_22_reset),
    .io_rd_valid(MemController_22_io_rd_valid),
    .io_wr_valid(MemController_22_io_wr_valid),
    .io_rd_data_valid(MemController_22_io_rd_data_valid),
    .io_rd_data_bits(MemController_22_io_rd_data_bits),
    .io_wr_data_valid(MemController_22_io_wr_data_valid),
    .io_wr_data_bits(MemController_22_io_wr_data_bits)
  );
  MemController_22 MemController_23 ( // @[pe.scala 303:15]
    .clock(MemController_23_clock),
    .reset(MemController_23_reset),
    .io_rd_valid(MemController_23_io_rd_valid),
    .io_wr_valid(MemController_23_io_wr_valid),
    .io_rd_data_valid(MemController_23_io_rd_data_valid),
    .io_rd_data_bits(MemController_23_io_rd_data_bits),
    .io_wr_data_valid(MemController_23_io_wr_data_valid),
    .io_wr_data_bits(MemController_23_io_wr_data_bits)
  );
  MemController_22 MemController_24 ( // @[pe.scala 303:15]
    .clock(MemController_24_clock),
    .reset(MemController_24_reset),
    .io_rd_valid(MemController_24_io_rd_valid),
    .io_wr_valid(MemController_24_io_wr_valid),
    .io_rd_data_valid(MemController_24_io_rd_data_valid),
    .io_rd_data_bits(MemController_24_io_rd_data_bits),
    .io_wr_data_valid(MemController_24_io_wr_data_valid),
    .io_wr_data_bits(MemController_24_io_wr_data_bits)
  );
  MemController_22 MemController_25 ( // @[pe.scala 303:15]
    .clock(MemController_25_clock),
    .reset(MemController_25_reset),
    .io_rd_valid(MemController_25_io_rd_valid),
    .io_wr_valid(MemController_25_io_wr_valid),
    .io_rd_data_valid(MemController_25_io_rd_data_valid),
    .io_rd_data_bits(MemController_25_io_rd_data_bits),
    .io_wr_data_valid(MemController_25_io_wr_data_valid),
    .io_wr_data_bits(MemController_25_io_wr_data_bits)
  );
  MemController_22 MemController_26 ( // @[pe.scala 303:15]
    .clock(MemController_26_clock),
    .reset(MemController_26_reset),
    .io_rd_valid(MemController_26_io_rd_valid),
    .io_wr_valid(MemController_26_io_wr_valid),
    .io_rd_data_valid(MemController_26_io_rd_data_valid),
    .io_rd_data_bits(MemController_26_io_rd_data_bits),
    .io_wr_data_valid(MemController_26_io_wr_data_valid),
    .io_wr_data_bits(MemController_26_io_wr_data_bits)
  );
  MemController_22 MemController_27 ( // @[pe.scala 303:15]
    .clock(MemController_27_clock),
    .reset(MemController_27_reset),
    .io_rd_valid(MemController_27_io_rd_valid),
    .io_wr_valid(MemController_27_io_wr_valid),
    .io_rd_data_valid(MemController_27_io_rd_data_valid),
    .io_rd_data_bits(MemController_27_io_rd_data_bits),
    .io_wr_data_valid(MemController_27_io_wr_data_valid),
    .io_wr_data_bits(MemController_27_io_wr_data_bits)
  );
  MemController_22 MemController_28 ( // @[pe.scala 303:15]
    .clock(MemController_28_clock),
    .reset(MemController_28_reset),
    .io_rd_valid(MemController_28_io_rd_valid),
    .io_wr_valid(MemController_28_io_wr_valid),
    .io_rd_data_valid(MemController_28_io_rd_data_valid),
    .io_rd_data_bits(MemController_28_io_rd_data_bits),
    .io_wr_data_valid(MemController_28_io_wr_data_valid),
    .io_wr_data_bits(MemController_28_io_wr_data_bits)
  );
  MemController_22 MemController_29 ( // @[pe.scala 303:15]
    .clock(MemController_29_clock),
    .reset(MemController_29_reset),
    .io_rd_valid(MemController_29_io_rd_valid),
    .io_wr_valid(MemController_29_io_wr_valid),
    .io_rd_data_valid(MemController_29_io_rd_data_valid),
    .io_rd_data_bits(MemController_29_io_rd_data_bits),
    .io_wr_data_valid(MemController_29_io_wr_data_valid),
    .io_wr_data_bits(MemController_29_io_wr_data_bits)
  );
  MemController_22 MemController_30 ( // @[pe.scala 303:15]
    .clock(MemController_30_clock),
    .reset(MemController_30_reset),
    .io_rd_valid(MemController_30_io_rd_valid),
    .io_wr_valid(MemController_30_io_wr_valid),
    .io_rd_data_valid(MemController_30_io_rd_data_valid),
    .io_rd_data_bits(MemController_30_io_rd_data_bits),
    .io_wr_data_valid(MemController_30_io_wr_data_valid),
    .io_wr_data_bits(MemController_30_io_wr_data_bits)
  );
  MemController_22 MemController_31 ( // @[pe.scala 303:15]
    .clock(MemController_31_clock),
    .reset(MemController_31_reset),
    .io_rd_valid(MemController_31_io_rd_valid),
    .io_wr_valid(MemController_31_io_wr_valid),
    .io_rd_data_valid(MemController_31_io_rd_data_valid),
    .io_rd_data_bits(MemController_31_io_rd_data_bits),
    .io_wr_data_valid(MemController_31_io_wr_data_valid),
    .io_wr_data_bits(MemController_31_io_wr_data_bits)
  );
  MemController_22 MemController_32 ( // @[pe.scala 303:15]
    .clock(MemController_32_clock),
    .reset(MemController_32_reset),
    .io_rd_valid(MemController_32_io_rd_valid),
    .io_wr_valid(MemController_32_io_wr_valid),
    .io_rd_data_valid(MemController_32_io_rd_data_valid),
    .io_rd_data_bits(MemController_32_io_rd_data_bits),
    .io_wr_data_valid(MemController_32_io_wr_data_valid),
    .io_wr_data_bits(MemController_32_io_wr_data_bits)
  );
  MemController_22 MemController_33 ( // @[pe.scala 303:15]
    .clock(MemController_33_clock),
    .reset(MemController_33_reset),
    .io_rd_valid(MemController_33_io_rd_valid),
    .io_wr_valid(MemController_33_io_wr_valid),
    .io_rd_data_valid(MemController_33_io_rd_data_valid),
    .io_rd_data_bits(MemController_33_io_rd_data_bits),
    .io_wr_data_valid(MemController_33_io_wr_data_valid),
    .io_wr_data_bits(MemController_33_io_wr_data_bits)
  );
  MemController_22 MemController_34 ( // @[pe.scala 303:15]
    .clock(MemController_34_clock),
    .reset(MemController_34_reset),
    .io_rd_valid(MemController_34_io_rd_valid),
    .io_wr_valid(MemController_34_io_wr_valid),
    .io_rd_data_valid(MemController_34_io_rd_data_valid),
    .io_rd_data_bits(MemController_34_io_rd_data_bits),
    .io_wr_data_valid(MemController_34_io_wr_data_valid),
    .io_wr_data_bits(MemController_34_io_wr_data_bits)
  );
  MemController_22 MemController_35 ( // @[pe.scala 303:15]
    .clock(MemController_35_clock),
    .reset(MemController_35_reset),
    .io_rd_valid(MemController_35_io_rd_valid),
    .io_wr_valid(MemController_35_io_wr_valid),
    .io_rd_data_valid(MemController_35_io_rd_data_valid),
    .io_rd_data_bits(MemController_35_io_rd_data_bits),
    .io_wr_data_valid(MemController_35_io_wr_data_valid),
    .io_wr_data_bits(MemController_35_io_wr_data_bits)
  );
  MemController_22 MemController_36 ( // @[pe.scala 303:15]
    .clock(MemController_36_clock),
    .reset(MemController_36_reset),
    .io_rd_valid(MemController_36_io_rd_valid),
    .io_wr_valid(MemController_36_io_wr_valid),
    .io_rd_data_valid(MemController_36_io_rd_data_valid),
    .io_rd_data_bits(MemController_36_io_rd_data_bits),
    .io_wr_data_valid(MemController_36_io_wr_data_valid),
    .io_wr_data_bits(MemController_36_io_wr_data_bits)
  );
  MemController_22 MemController_37 ( // @[pe.scala 303:15]
    .clock(MemController_37_clock),
    .reset(MemController_37_reset),
    .io_rd_valid(MemController_37_io_rd_valid),
    .io_wr_valid(MemController_37_io_wr_valid),
    .io_rd_data_valid(MemController_37_io_rd_data_valid),
    .io_rd_data_bits(MemController_37_io_rd_data_bits),
    .io_wr_data_valid(MemController_37_io_wr_data_valid),
    .io_wr_data_bits(MemController_37_io_wr_data_bits)
  );
  MemController_22 MemController_38 ( // @[pe.scala 303:15]
    .clock(MemController_38_clock),
    .reset(MemController_38_reset),
    .io_rd_valid(MemController_38_io_rd_valid),
    .io_wr_valid(MemController_38_io_wr_valid),
    .io_rd_data_valid(MemController_38_io_rd_data_valid),
    .io_rd_data_bits(MemController_38_io_rd_data_bits),
    .io_wr_data_valid(MemController_38_io_wr_data_valid),
    .io_wr_data_bits(MemController_38_io_wr_data_bits)
  );
  MemController_22 MemController_39 ( // @[pe.scala 303:15]
    .clock(MemController_39_clock),
    .reset(MemController_39_reset),
    .io_rd_valid(MemController_39_io_rd_valid),
    .io_wr_valid(MemController_39_io_wr_valid),
    .io_rd_data_valid(MemController_39_io_rd_data_valid),
    .io_rd_data_bits(MemController_39_io_rd_data_bits),
    .io_wr_data_valid(MemController_39_io_wr_data_valid),
    .io_wr_data_bits(MemController_39_io_wr_data_bits)
  );
  MemController_22 MemController_40 ( // @[pe.scala 303:15]
    .clock(MemController_40_clock),
    .reset(MemController_40_reset),
    .io_rd_valid(MemController_40_io_rd_valid),
    .io_wr_valid(MemController_40_io_wr_valid),
    .io_rd_data_valid(MemController_40_io_rd_data_valid),
    .io_rd_data_bits(MemController_40_io_rd_data_bits),
    .io_wr_data_valid(MemController_40_io_wr_data_valid),
    .io_wr_data_bits(MemController_40_io_wr_data_bits)
  );
  MemController_22 MemController_41 ( // @[pe.scala 303:15]
    .clock(MemController_41_clock),
    .reset(MemController_41_reset),
    .io_rd_valid(MemController_41_io_rd_valid),
    .io_wr_valid(MemController_41_io_wr_valid),
    .io_rd_data_valid(MemController_41_io_rd_data_valid),
    .io_rd_data_bits(MemController_41_io_rd_data_bits),
    .io_wr_data_valid(MemController_41_io_wr_data_valid),
    .io_wr_data_bits(MemController_41_io_wr_data_bits)
  );
  MemController_22 MemController_42 ( // @[pe.scala 303:15]
    .clock(MemController_42_clock),
    .reset(MemController_42_reset),
    .io_rd_valid(MemController_42_io_rd_valid),
    .io_wr_valid(MemController_42_io_wr_valid),
    .io_rd_data_valid(MemController_42_io_rd_data_valid),
    .io_rd_data_bits(MemController_42_io_rd_data_bits),
    .io_wr_data_valid(MemController_42_io_wr_data_valid),
    .io_wr_data_bits(MemController_42_io_wr_data_bits)
  );
  MemController_22 MemController_43 ( // @[pe.scala 303:15]
    .clock(MemController_43_clock),
    .reset(MemController_43_reset),
    .io_rd_valid(MemController_43_io_rd_valid),
    .io_wr_valid(MemController_43_io_wr_valid),
    .io_rd_data_valid(MemController_43_io_rd_data_valid),
    .io_rd_data_bits(MemController_43_io_rd_data_bits),
    .io_wr_data_valid(MemController_43_io_wr_data_valid),
    .io_wr_data_bits(MemController_43_io_wr_data_bits)
  );
  MemController_22 MemController_44 ( // @[pe.scala 303:15]
    .clock(MemController_44_clock),
    .reset(MemController_44_reset),
    .io_rd_valid(MemController_44_io_rd_valid),
    .io_wr_valid(MemController_44_io_wr_valid),
    .io_rd_data_valid(MemController_44_io_rd_data_valid),
    .io_rd_data_bits(MemController_44_io_rd_data_bits),
    .io_wr_data_valid(MemController_44_io_wr_data_valid),
    .io_wr_data_bits(MemController_44_io_wr_data_bits)
  );
  MemController_22 MemController_45 ( // @[pe.scala 303:15]
    .clock(MemController_45_clock),
    .reset(MemController_45_reset),
    .io_rd_valid(MemController_45_io_rd_valid),
    .io_wr_valid(MemController_45_io_wr_valid),
    .io_rd_data_valid(MemController_45_io_rd_data_valid),
    .io_rd_data_bits(MemController_45_io_rd_data_bits),
    .io_wr_data_valid(MemController_45_io_wr_data_valid),
    .io_wr_data_bits(MemController_45_io_wr_data_bits)
  );
  MemController_22 MemController_46 ( // @[pe.scala 303:15]
    .clock(MemController_46_clock),
    .reset(MemController_46_reset),
    .io_rd_valid(MemController_46_io_rd_valid),
    .io_wr_valid(MemController_46_io_wr_valid),
    .io_rd_data_valid(MemController_46_io_rd_data_valid),
    .io_rd_data_bits(MemController_46_io_rd_data_bits),
    .io_wr_data_valid(MemController_46_io_wr_data_valid),
    .io_wr_data_bits(MemController_46_io_wr_data_bits)
  );
  MemController_22 MemController_47 ( // @[pe.scala 303:15]
    .clock(MemController_47_clock),
    .reset(MemController_47_reset),
    .io_rd_valid(MemController_47_io_rd_valid),
    .io_wr_valid(MemController_47_io_wr_valid),
    .io_rd_data_valid(MemController_47_io_rd_data_valid),
    .io_rd_data_bits(MemController_47_io_rd_data_bits),
    .io_wr_data_valid(MemController_47_io_wr_data_valid),
    .io_wr_data_bits(MemController_47_io_wr_data_bits)
  );
  MemController_22 MemController_48 ( // @[pe.scala 303:15]
    .clock(MemController_48_clock),
    .reset(MemController_48_reset),
    .io_rd_valid(MemController_48_io_rd_valid),
    .io_wr_valid(MemController_48_io_wr_valid),
    .io_rd_data_valid(MemController_48_io_rd_data_valid),
    .io_rd_data_bits(MemController_48_io_rd_data_bits),
    .io_wr_data_valid(MemController_48_io_wr_data_valid),
    .io_wr_data_bits(MemController_48_io_wr_data_bits)
  );
  MemController_22 MemController_49 ( // @[pe.scala 303:15]
    .clock(MemController_49_clock),
    .reset(MemController_49_reset),
    .io_rd_valid(MemController_49_io_rd_valid),
    .io_wr_valid(MemController_49_io_wr_valid),
    .io_rd_data_valid(MemController_49_io_rd_data_valid),
    .io_rd_data_bits(MemController_49_io_rd_data_bits),
    .io_wr_data_valid(MemController_49_io_wr_data_valid),
    .io_wr_data_bits(MemController_49_io_wr_data_bits)
  );
  MemController_22 MemController_50 ( // @[pe.scala 303:15]
    .clock(MemController_50_clock),
    .reset(MemController_50_reset),
    .io_rd_valid(MemController_50_io_rd_valid),
    .io_wr_valid(MemController_50_io_wr_valid),
    .io_rd_data_valid(MemController_50_io_rd_data_valid),
    .io_rd_data_bits(MemController_50_io_rd_data_bits),
    .io_wr_data_valid(MemController_50_io_wr_data_valid),
    .io_wr_data_bits(MemController_50_io_wr_data_bits)
  );
  MemController_22 MemController_51 ( // @[pe.scala 303:15]
    .clock(MemController_51_clock),
    .reset(MemController_51_reset),
    .io_rd_valid(MemController_51_io_rd_valid),
    .io_wr_valid(MemController_51_io_wr_valid),
    .io_rd_data_valid(MemController_51_io_rd_data_valid),
    .io_rd_data_bits(MemController_51_io_rd_data_bits),
    .io_wr_data_valid(MemController_51_io_wr_data_valid),
    .io_wr_data_bits(MemController_51_io_wr_data_bits)
  );
  MemController_52 MemController_52 ( // @[pe.scala 301:15]
    .clock(MemController_52_clock),
    .reset(MemController_52_reset),
    .io_rd_valid(MemController_52_io_rd_valid),
    .io_wr_valid(MemController_52_io_wr_valid),
    .io_rd_data_valid(MemController_52_io_rd_data_valid),
    .io_rd_data_bits(MemController_52_io_rd_data_bits),
    .io_wr_data_valid(MemController_52_io_wr_data_valid),
    .io_wr_data_bits(MemController_52_io_wr_data_bits)
  );
  MemController_52 MemController_53 ( // @[pe.scala 301:15]
    .clock(MemController_53_clock),
    .reset(MemController_53_reset),
    .io_rd_valid(MemController_53_io_rd_valid),
    .io_wr_valid(MemController_53_io_wr_valid),
    .io_rd_data_valid(MemController_53_io_rd_data_valid),
    .io_rd_data_bits(MemController_53_io_rd_data_bits),
    .io_wr_data_valid(MemController_53_io_wr_data_valid),
    .io_wr_data_bits(MemController_53_io_wr_data_bits)
  );
  MemController_52 MemController_54 ( // @[pe.scala 301:15]
    .clock(MemController_54_clock),
    .reset(MemController_54_reset),
    .io_rd_valid(MemController_54_io_rd_valid),
    .io_wr_valid(MemController_54_io_wr_valid),
    .io_rd_data_valid(MemController_54_io_rd_data_valid),
    .io_rd_data_bits(MemController_54_io_rd_data_bits),
    .io_wr_data_valid(MemController_54_io_wr_data_valid),
    .io_wr_data_bits(MemController_54_io_wr_data_bits)
  );
  MemController_52 MemController_55 ( // @[pe.scala 301:15]
    .clock(MemController_55_clock),
    .reset(MemController_55_reset),
    .io_rd_valid(MemController_55_io_rd_valid),
    .io_wr_valid(MemController_55_io_wr_valid),
    .io_rd_data_valid(MemController_55_io_rd_data_valid),
    .io_rd_data_bits(MemController_55_io_rd_data_bits),
    .io_wr_data_valid(MemController_55_io_wr_data_valid),
    .io_wr_data_bits(MemController_55_io_wr_data_bits)
  );
  MemController_52 MemController_56 ( // @[pe.scala 301:15]
    .clock(MemController_56_clock),
    .reset(MemController_56_reset),
    .io_rd_valid(MemController_56_io_rd_valid),
    .io_wr_valid(MemController_56_io_wr_valid),
    .io_rd_data_valid(MemController_56_io_rd_data_valid),
    .io_rd_data_bits(MemController_56_io_rd_data_bits),
    .io_wr_data_valid(MemController_56_io_wr_data_valid),
    .io_wr_data_bits(MemController_56_io_wr_data_bits)
  );
  MemController_52 MemController_57 ( // @[pe.scala 301:15]
    .clock(MemController_57_clock),
    .reset(MemController_57_reset),
    .io_rd_valid(MemController_57_io_rd_valid),
    .io_wr_valid(MemController_57_io_wr_valid),
    .io_rd_data_valid(MemController_57_io_rd_data_valid),
    .io_rd_data_bits(MemController_57_io_rd_data_bits),
    .io_wr_data_valid(MemController_57_io_wr_data_valid),
    .io_wr_data_bits(MemController_57_io_wr_data_bits)
  );
  MemController_52 MemController_58 ( // @[pe.scala 301:15]
    .clock(MemController_58_clock),
    .reset(MemController_58_reset),
    .io_rd_valid(MemController_58_io_rd_valid),
    .io_wr_valid(MemController_58_io_wr_valid),
    .io_rd_data_valid(MemController_58_io_rd_data_valid),
    .io_rd_data_bits(MemController_58_io_rd_data_bits),
    .io_wr_data_valid(MemController_58_io_wr_data_valid),
    .io_wr_data_bits(MemController_58_io_wr_data_bits)
  );
  MemController_52 MemController_59 ( // @[pe.scala 301:15]
    .clock(MemController_59_clock),
    .reset(MemController_59_reset),
    .io_rd_valid(MemController_59_io_rd_valid),
    .io_wr_valid(MemController_59_io_wr_valid),
    .io_rd_data_valid(MemController_59_io_rd_data_valid),
    .io_rd_data_bits(MemController_59_io_rd_data_bits),
    .io_wr_data_valid(MemController_59_io_wr_data_valid),
    .io_wr_data_bits(MemController_59_io_wr_data_bits)
  );
  MemController_52 MemController_60 ( // @[pe.scala 301:15]
    .clock(MemController_60_clock),
    .reset(MemController_60_reset),
    .io_rd_valid(MemController_60_io_rd_valid),
    .io_wr_valid(MemController_60_io_wr_valid),
    .io_rd_data_valid(MemController_60_io_rd_data_valid),
    .io_rd_data_bits(MemController_60_io_rd_data_bits),
    .io_wr_data_valid(MemController_60_io_wr_data_valid),
    .io_wr_data_bits(MemController_60_io_wr_data_bits)
  );
  MemController_52 MemController_61 ( // @[pe.scala 301:15]
    .clock(MemController_61_clock),
    .reset(MemController_61_reset),
    .io_rd_valid(MemController_61_io_rd_valid),
    .io_wr_valid(MemController_61_io_wr_valid),
    .io_rd_data_valid(MemController_61_io_rd_data_valid),
    .io_rd_data_bits(MemController_61_io_rd_data_bits),
    .io_wr_data_valid(MemController_61_io_wr_data_valid),
    .io_wr_data_bits(MemController_61_io_wr_data_bits)
  );
  MemController_52 MemController_62 ( // @[pe.scala 301:15]
    .clock(MemController_62_clock),
    .reset(MemController_62_reset),
    .io_rd_valid(MemController_62_io_rd_valid),
    .io_wr_valid(MemController_62_io_wr_valid),
    .io_rd_data_valid(MemController_62_io_rd_data_valid),
    .io_rd_data_bits(MemController_62_io_rd_data_bits),
    .io_wr_data_valid(MemController_62_io_wr_data_valid),
    .io_wr_data_bits(MemController_62_io_wr_data_bits)
  );
  MemController_52 MemController_63 ( // @[pe.scala 301:15]
    .clock(MemController_63_clock),
    .reset(MemController_63_reset),
    .io_rd_valid(MemController_63_io_rd_valid),
    .io_wr_valid(MemController_63_io_wr_valid),
    .io_rd_data_valid(MemController_63_io_rd_data_valid),
    .io_rd_data_bits(MemController_63_io_rd_data_bits),
    .io_wr_data_valid(MemController_63_io_wr_data_valid),
    .io_wr_data_bits(MemController_63_io_wr_data_bits)
  );
  MemController_52 MemController_64 ( // @[pe.scala 301:15]
    .clock(MemController_64_clock),
    .reset(MemController_64_reset),
    .io_rd_valid(MemController_64_io_rd_valid),
    .io_wr_valid(MemController_64_io_wr_valid),
    .io_rd_data_valid(MemController_64_io_rd_data_valid),
    .io_rd_data_bits(MemController_64_io_rd_data_bits),
    .io_wr_data_valid(MemController_64_io_wr_data_valid),
    .io_wr_data_bits(MemController_64_io_wr_data_bits)
  );
  MemController_52 MemController_65 ( // @[pe.scala 301:15]
    .clock(MemController_65_clock),
    .reset(MemController_65_reset),
    .io_rd_valid(MemController_65_io_rd_valid),
    .io_wr_valid(MemController_65_io_wr_valid),
    .io_rd_data_valid(MemController_65_io_rd_data_valid),
    .io_rd_data_bits(MemController_65_io_rd_data_bits),
    .io_wr_data_valid(MemController_65_io_wr_data_valid),
    .io_wr_data_bits(MemController_65_io_wr_data_bits)
  );
  MemController_52 MemController_66 ( // @[pe.scala 301:15]
    .clock(MemController_66_clock),
    .reset(MemController_66_reset),
    .io_rd_valid(MemController_66_io_rd_valid),
    .io_wr_valid(MemController_66_io_wr_valid),
    .io_rd_data_valid(MemController_66_io_rd_data_valid),
    .io_rd_data_bits(MemController_66_io_rd_data_bits),
    .io_wr_data_valid(MemController_66_io_wr_data_valid),
    .io_wr_data_bits(MemController_66_io_wr_data_bits)
  );
  MemController_52 MemController_67 ( // @[pe.scala 301:15]
    .clock(MemController_67_clock),
    .reset(MemController_67_reset),
    .io_rd_valid(MemController_67_io_rd_valid),
    .io_wr_valid(MemController_67_io_wr_valid),
    .io_rd_data_valid(MemController_67_io_rd_data_valid),
    .io_rd_data_bits(MemController_67_io_rd_data_bits),
    .io_wr_data_valid(MemController_67_io_wr_data_valid),
    .io_wr_data_bits(MemController_67_io_wr_data_bits)
  );
  MemController_52 MemController_68 ( // @[pe.scala 301:15]
    .clock(MemController_68_clock),
    .reset(MemController_68_reset),
    .io_rd_valid(MemController_68_io_rd_valid),
    .io_wr_valid(MemController_68_io_wr_valid),
    .io_rd_data_valid(MemController_68_io_rd_data_valid),
    .io_rd_data_bits(MemController_68_io_rd_data_bits),
    .io_wr_data_valid(MemController_68_io_wr_data_valid),
    .io_wr_data_bits(MemController_68_io_wr_data_bits)
  );
  MemController_52 MemController_69 ( // @[pe.scala 301:15]
    .clock(MemController_69_clock),
    .reset(MemController_69_reset),
    .io_rd_valid(MemController_69_io_rd_valid),
    .io_wr_valid(MemController_69_io_wr_valid),
    .io_rd_data_valid(MemController_69_io_rd_data_valid),
    .io_rd_data_bits(MemController_69_io_rd_data_bits),
    .io_wr_data_valid(MemController_69_io_wr_data_valid),
    .io_wr_data_bits(MemController_69_io_wr_data_bits)
  );
  MemController_52 MemController_70 ( // @[pe.scala 301:15]
    .clock(MemController_70_clock),
    .reset(MemController_70_reset),
    .io_rd_valid(MemController_70_io_rd_valid),
    .io_wr_valid(MemController_70_io_wr_valid),
    .io_rd_data_valid(MemController_70_io_rd_data_valid),
    .io_rd_data_bits(MemController_70_io_rd_data_bits),
    .io_wr_data_valid(MemController_70_io_wr_data_valid),
    .io_wr_data_bits(MemController_70_io_wr_data_bits)
  );
  MemController_52 MemController_71 ( // @[pe.scala 301:15]
    .clock(MemController_71_clock),
    .reset(MemController_71_reset),
    .io_rd_valid(MemController_71_io_rd_valid),
    .io_wr_valid(MemController_71_io_wr_valid),
    .io_rd_data_valid(MemController_71_io_rd_data_valid),
    .io_rd_data_bits(MemController_71_io_rd_data_bits),
    .io_wr_data_valid(MemController_71_io_wr_data_valid),
    .io_wr_data_bits(MemController_71_io_wr_data_bits)
  );
  MemController_52 MemController_72 ( // @[pe.scala 301:15]
    .clock(MemController_72_clock),
    .reset(MemController_72_reset),
    .io_rd_valid(MemController_72_io_rd_valid),
    .io_wr_valid(MemController_72_io_wr_valid),
    .io_rd_data_valid(MemController_72_io_rd_data_valid),
    .io_rd_data_bits(MemController_72_io_rd_data_bits),
    .io_wr_data_valid(MemController_72_io_wr_data_valid),
    .io_wr_data_bits(MemController_72_io_wr_data_bits)
  );
  MemController_52 MemController_73 ( // @[pe.scala 301:15]
    .clock(MemController_73_clock),
    .reset(MemController_73_reset),
    .io_rd_valid(MemController_73_io_rd_valid),
    .io_wr_valid(MemController_73_io_wr_valid),
    .io_rd_data_valid(MemController_73_io_rd_data_valid),
    .io_rd_data_bits(MemController_73_io_rd_data_bits),
    .io_wr_data_valid(MemController_73_io_wr_data_valid),
    .io_wr_data_bits(MemController_73_io_wr_data_bits)
  );
  MemController_52 MemController_74 ( // @[pe.scala 301:15]
    .clock(MemController_74_clock),
    .reset(MemController_74_reset),
    .io_rd_valid(MemController_74_io_rd_valid),
    .io_wr_valid(MemController_74_io_wr_valid),
    .io_rd_data_valid(MemController_74_io_rd_data_valid),
    .io_rd_data_bits(MemController_74_io_rd_data_bits),
    .io_wr_data_valid(MemController_74_io_wr_data_valid),
    .io_wr_data_bits(MemController_74_io_wr_data_bits)
  );
  MemController_52 MemController_75 ( // @[pe.scala 301:15]
    .clock(MemController_75_clock),
    .reset(MemController_75_reset),
    .io_rd_valid(MemController_75_io_rd_valid),
    .io_wr_valid(MemController_75_io_wr_valid),
    .io_rd_data_valid(MemController_75_io_rd_data_valid),
    .io_rd_data_bits(MemController_75_io_rd_data_bits),
    .io_wr_data_valid(MemController_75_io_wr_data_valid),
    .io_wr_data_bits(MemController_75_io_wr_data_bits)
  );
  MemController_52 MemController_76 ( // @[pe.scala 301:15]
    .clock(MemController_76_clock),
    .reset(MemController_76_reset),
    .io_rd_valid(MemController_76_io_rd_valid),
    .io_wr_valid(MemController_76_io_wr_valid),
    .io_rd_data_valid(MemController_76_io_rd_data_valid),
    .io_rd_data_bits(MemController_76_io_rd_data_bits),
    .io_wr_data_valid(MemController_76_io_wr_data_valid),
    .io_wr_data_bits(MemController_76_io_wr_data_bits)
  );
  MemController_52 MemController_77 ( // @[pe.scala 301:15]
    .clock(MemController_77_clock),
    .reset(MemController_77_reset),
    .io_rd_valid(MemController_77_io_rd_valid),
    .io_wr_valid(MemController_77_io_wr_valid),
    .io_rd_data_valid(MemController_77_io_rd_data_valid),
    .io_rd_data_bits(MemController_77_io_rd_data_bits),
    .io_wr_data_valid(MemController_77_io_wr_data_valid),
    .io_wr_data_bits(MemController_77_io_wr_data_bits)
  );
  MemController_52 MemController_78 ( // @[pe.scala 301:15]
    .clock(MemController_78_clock),
    .reset(MemController_78_reset),
    .io_rd_valid(MemController_78_io_rd_valid),
    .io_wr_valid(MemController_78_io_wr_valid),
    .io_rd_data_valid(MemController_78_io_rd_data_valid),
    .io_rd_data_bits(MemController_78_io_rd_data_bits),
    .io_wr_data_valid(MemController_78_io_wr_data_valid),
    .io_wr_data_bits(MemController_78_io_wr_data_bits)
  );
  MemController_52 MemController_79 ( // @[pe.scala 301:15]
    .clock(MemController_79_clock),
    .reset(MemController_79_reset),
    .io_rd_valid(MemController_79_io_rd_valid),
    .io_wr_valid(MemController_79_io_wr_valid),
    .io_rd_data_valid(MemController_79_io_rd_data_valid),
    .io_rd_data_bits(MemController_79_io_rd_data_bits),
    .io_wr_data_valid(MemController_79_io_wr_data_valid),
    .io_wr_data_bits(MemController_79_io_wr_data_bits)
  );
  MemController_52 MemController_80 ( // @[pe.scala 301:15]
    .clock(MemController_80_clock),
    .reset(MemController_80_reset),
    .io_rd_valid(MemController_80_io_rd_valid),
    .io_wr_valid(MemController_80_io_wr_valid),
    .io_rd_data_valid(MemController_80_io_rd_data_valid),
    .io_rd_data_bits(MemController_80_io_rd_data_bits),
    .io_wr_data_valid(MemController_80_io_wr_data_valid),
    .io_wr_data_bits(MemController_80_io_wr_data_bits)
  );
  MemController_52 MemController_81 ( // @[pe.scala 301:15]
    .clock(MemController_81_clock),
    .reset(MemController_81_reset),
    .io_rd_valid(MemController_81_io_rd_valid),
    .io_wr_valid(MemController_81_io_wr_valid),
    .io_rd_data_valid(MemController_81_io_rd_data_valid),
    .io_rd_data_bits(MemController_81_io_rd_data_bits),
    .io_wr_data_valid(MemController_81_io_wr_data_valid),
    .io_wr_data_bits(MemController_81_io_wr_data_bits)
  );
  assign io_data_2_out_0_valid = MemController_52_io_rd_data_valid; // @[pe.scala 318:31]
  assign io_data_2_out_0_bits = MemController_52_io_rd_data_bits; // @[pe.scala 318:31]
  assign io_data_2_out_1_valid = MemController_53_io_rd_data_valid; // @[pe.scala 318:31]
  assign io_data_2_out_1_bits = MemController_53_io_rd_data_bits; // @[pe.scala 318:31]
  assign io_data_2_out_2_valid = MemController_54_io_rd_data_valid; // @[pe.scala 318:31]
  assign io_data_2_out_2_bits = MemController_54_io_rd_data_bits; // @[pe.scala 318:31]
  assign io_data_2_out_3_valid = MemController_55_io_rd_data_valid; // @[pe.scala 318:31]
  assign io_data_2_out_3_bits = MemController_55_io_rd_data_bits; // @[pe.scala 318:31]
  assign io_data_2_out_4_valid = MemController_56_io_rd_data_valid; // @[pe.scala 318:31]
  assign io_data_2_out_4_bits = MemController_56_io_rd_data_bits; // @[pe.scala 318:31]
  assign io_data_2_out_5_valid = MemController_57_io_rd_data_valid; // @[pe.scala 318:31]
  assign io_data_2_out_5_bits = MemController_57_io_rd_data_bits; // @[pe.scala 318:31]
  assign io_data_2_out_6_valid = MemController_58_io_rd_data_valid; // @[pe.scala 318:31]
  assign io_data_2_out_6_bits = MemController_58_io_rd_data_bits; // @[pe.scala 318:31]
  assign io_data_2_out_7_valid = MemController_59_io_rd_data_valid; // @[pe.scala 318:31]
  assign io_data_2_out_7_bits = MemController_59_io_rd_data_bits; // @[pe.scala 318:31]
  assign io_data_2_out_8_valid = MemController_60_io_rd_data_valid; // @[pe.scala 318:31]
  assign io_data_2_out_8_bits = MemController_60_io_rd_data_bits; // @[pe.scala 318:31]
  assign io_data_2_out_9_valid = MemController_61_io_rd_data_valid; // @[pe.scala 318:31]
  assign io_data_2_out_9_bits = MemController_61_io_rd_data_bits; // @[pe.scala 318:31]
  assign io_data_2_out_10_valid = MemController_62_io_rd_data_valid; // @[pe.scala 318:31]
  assign io_data_2_out_10_bits = MemController_62_io_rd_data_bits; // @[pe.scala 318:31]
  assign io_data_2_out_11_valid = MemController_63_io_rd_data_valid; // @[pe.scala 318:31]
  assign io_data_2_out_11_bits = MemController_63_io_rd_data_bits; // @[pe.scala 318:31]
  assign io_data_2_out_12_valid = MemController_64_io_rd_data_valid; // @[pe.scala 318:31]
  assign io_data_2_out_12_bits = MemController_64_io_rd_data_bits; // @[pe.scala 318:31]
  assign io_data_2_out_13_valid = MemController_65_io_rd_data_valid; // @[pe.scala 318:31]
  assign io_data_2_out_13_bits = MemController_65_io_rd_data_bits; // @[pe.scala 318:31]
  assign io_data_2_out_14_valid = MemController_66_io_rd_data_valid; // @[pe.scala 318:31]
  assign io_data_2_out_14_bits = MemController_66_io_rd_data_bits; // @[pe.scala 318:31]
  assign io_data_2_out_15_valid = MemController_67_io_rd_data_valid; // @[pe.scala 318:31]
  assign io_data_2_out_15_bits = MemController_67_io_rd_data_bits; // @[pe.scala 318:31]
  assign io_data_2_out_16_valid = MemController_68_io_rd_data_valid; // @[pe.scala 318:31]
  assign io_data_2_out_16_bits = MemController_68_io_rd_data_bits; // @[pe.scala 318:31]
  assign io_data_2_out_17_valid = MemController_69_io_rd_data_valid; // @[pe.scala 318:31]
  assign io_data_2_out_17_bits = MemController_69_io_rd_data_bits; // @[pe.scala 318:31]
  assign io_data_2_out_18_valid = MemController_70_io_rd_data_valid; // @[pe.scala 318:31]
  assign io_data_2_out_18_bits = MemController_70_io_rd_data_bits; // @[pe.scala 318:31]
  assign io_data_2_out_19_valid = MemController_71_io_rd_data_valid; // @[pe.scala 318:31]
  assign io_data_2_out_19_bits = MemController_71_io_rd_data_bits; // @[pe.scala 318:31]
  assign io_data_2_out_20_valid = MemController_72_io_rd_data_valid; // @[pe.scala 318:31]
  assign io_data_2_out_20_bits = MemController_72_io_rd_data_bits; // @[pe.scala 318:31]
  assign io_data_2_out_21_valid = MemController_73_io_rd_data_valid; // @[pe.scala 318:31]
  assign io_data_2_out_21_bits = MemController_73_io_rd_data_bits; // @[pe.scala 318:31]
  assign io_data_2_out_22_valid = MemController_74_io_rd_data_valid; // @[pe.scala 318:31]
  assign io_data_2_out_22_bits = MemController_74_io_rd_data_bits; // @[pe.scala 318:31]
  assign io_data_2_out_23_valid = MemController_75_io_rd_data_valid; // @[pe.scala 318:31]
  assign io_data_2_out_23_bits = MemController_75_io_rd_data_bits; // @[pe.scala 318:31]
  assign io_data_2_out_24_valid = MemController_76_io_rd_data_valid; // @[pe.scala 318:31]
  assign io_data_2_out_24_bits = MemController_76_io_rd_data_bits; // @[pe.scala 318:31]
  assign io_data_2_out_25_valid = MemController_77_io_rd_data_valid; // @[pe.scala 318:31]
  assign io_data_2_out_25_bits = MemController_77_io_rd_data_bits; // @[pe.scala 318:31]
  assign io_data_2_out_26_valid = MemController_78_io_rd_data_valid; // @[pe.scala 318:31]
  assign io_data_2_out_26_bits = MemController_78_io_rd_data_bits; // @[pe.scala 318:31]
  assign io_data_2_out_27_valid = MemController_79_io_rd_data_valid; // @[pe.scala 318:31]
  assign io_data_2_out_27_bits = MemController_79_io_rd_data_bits; // @[pe.scala 318:31]
  assign io_data_2_out_28_valid = MemController_80_io_rd_data_valid; // @[pe.scala 318:31]
  assign io_data_2_out_28_bits = MemController_80_io_rd_data_bits; // @[pe.scala 318:31]
  assign io_data_2_out_29_valid = MemController_81_io_rd_data_valid; // @[pe.scala 318:31]
  assign io_data_2_out_29_bits = MemController_81_io_rd_data_bits; // @[pe.scala 318:31]
  assign MultiDimTime_clock = clock;
  assign MultiDimTime_reset = reset;
  assign MultiDimTime_io_in = io_exec_valid; // @[pe.scala 257:16]
  assign PE_clock = clock;
  assign PE_reset = reset;
  assign PE_io_data_2_sig_stat2trans = PENetwork_52_io_to_pes_0_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_io_data_1_in_valid = PENetwork_22_io_to_pes_0_in_valid; // @[pe.scala 264:34]
  assign PE_io_data_1_in_bits = PENetwork_22_io_to_pes_0_in_bits; // @[pe.scala 264:34]
  assign PE_io_data_0_in_valid = PENetwork_io_to_pes_0_in_valid; // @[pe.scala 264:34]
  assign PE_io_data_0_in_bits = PENetwork_io_to_pes_0_in_bits; // @[pe.scala 264:34]
  assign PE_1_clock = clock;
  assign PE_1_reset = reset;
  assign PE_1_io_data_2_sig_stat2trans = PENetwork_52_io_to_pes_1_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_1_io_data_1_in_valid = PENetwork_22_io_to_pes_1_in_valid; // @[pe.scala 264:34]
  assign PE_1_io_data_1_in_bits = PENetwork_22_io_to_pes_1_in_bits; // @[pe.scala 264:34]
  assign PE_1_io_data_0_in_valid = PENetwork_1_io_to_pes_0_in_valid; // @[pe.scala 264:34]
  assign PE_1_io_data_0_in_bits = PENetwork_1_io_to_pes_0_in_bits; // @[pe.scala 264:34]
  assign PE_2_clock = clock;
  assign PE_2_reset = reset;
  assign PE_2_io_data_2_sig_stat2trans = PENetwork_52_io_to_pes_2_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_2_io_data_1_in_valid = PENetwork_22_io_to_pes_2_in_valid; // @[pe.scala 264:34]
  assign PE_2_io_data_1_in_bits = PENetwork_22_io_to_pes_2_in_bits; // @[pe.scala 264:34]
  assign PE_2_io_data_0_in_valid = PENetwork_2_io_to_pes_0_in_valid; // @[pe.scala 264:34]
  assign PE_2_io_data_0_in_bits = PENetwork_2_io_to_pes_0_in_bits; // @[pe.scala 264:34]
  assign PE_3_clock = clock;
  assign PE_3_reset = reset;
  assign PE_3_io_data_2_sig_stat2trans = PENetwork_52_io_to_pes_3_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_3_io_data_1_in_valid = PENetwork_22_io_to_pes_3_in_valid; // @[pe.scala 264:34]
  assign PE_3_io_data_1_in_bits = PENetwork_22_io_to_pes_3_in_bits; // @[pe.scala 264:34]
  assign PE_3_io_data_0_in_valid = PENetwork_3_io_to_pes_0_in_valid; // @[pe.scala 264:34]
  assign PE_3_io_data_0_in_bits = PENetwork_3_io_to_pes_0_in_bits; // @[pe.scala 264:34]
  assign PE_4_clock = clock;
  assign PE_4_reset = reset;
  assign PE_4_io_data_2_sig_stat2trans = PENetwork_52_io_to_pes_4_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_4_io_data_1_in_valid = PENetwork_22_io_to_pes_4_in_valid; // @[pe.scala 264:34]
  assign PE_4_io_data_1_in_bits = PENetwork_22_io_to_pes_4_in_bits; // @[pe.scala 264:34]
  assign PE_4_io_data_0_in_valid = PENetwork_4_io_to_pes_0_in_valid; // @[pe.scala 264:34]
  assign PE_4_io_data_0_in_bits = PENetwork_4_io_to_pes_0_in_bits; // @[pe.scala 264:34]
  assign PE_5_clock = clock;
  assign PE_5_reset = reset;
  assign PE_5_io_data_2_sig_stat2trans = PENetwork_52_io_to_pes_5_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_5_io_data_1_in_valid = PENetwork_22_io_to_pes_5_in_valid; // @[pe.scala 264:34]
  assign PE_5_io_data_1_in_bits = PENetwork_22_io_to_pes_5_in_bits; // @[pe.scala 264:34]
  assign PE_5_io_data_0_in_valid = PENetwork_5_io_to_pes_0_in_valid; // @[pe.scala 264:34]
  assign PE_5_io_data_0_in_bits = PENetwork_5_io_to_pes_0_in_bits; // @[pe.scala 264:34]
  assign PE_6_clock = clock;
  assign PE_6_reset = reset;
  assign PE_6_io_data_2_sig_stat2trans = PENetwork_52_io_to_pes_6_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_6_io_data_1_in_valid = PENetwork_22_io_to_pes_6_in_valid; // @[pe.scala 264:34]
  assign PE_6_io_data_1_in_bits = PENetwork_22_io_to_pes_6_in_bits; // @[pe.scala 264:34]
  assign PE_6_io_data_0_in_valid = PENetwork_6_io_to_pes_0_in_valid; // @[pe.scala 264:34]
  assign PE_6_io_data_0_in_bits = PENetwork_6_io_to_pes_0_in_bits; // @[pe.scala 264:34]
  assign PE_7_clock = clock;
  assign PE_7_reset = reset;
  assign PE_7_io_data_2_sig_stat2trans = PENetwork_52_io_to_pes_7_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_7_io_data_1_in_valid = PENetwork_22_io_to_pes_7_in_valid; // @[pe.scala 264:34]
  assign PE_7_io_data_1_in_bits = PENetwork_22_io_to_pes_7_in_bits; // @[pe.scala 264:34]
  assign PE_7_io_data_0_in_valid = PENetwork_7_io_to_pes_0_in_valid; // @[pe.scala 264:34]
  assign PE_7_io_data_0_in_bits = PENetwork_7_io_to_pes_0_in_bits; // @[pe.scala 264:34]
  assign PE_8_clock = clock;
  assign PE_8_reset = reset;
  assign PE_8_io_data_2_sig_stat2trans = PENetwork_52_io_to_pes_8_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_8_io_data_1_in_valid = PENetwork_22_io_to_pes_8_in_valid; // @[pe.scala 264:34]
  assign PE_8_io_data_1_in_bits = PENetwork_22_io_to_pes_8_in_bits; // @[pe.scala 264:34]
  assign PE_8_io_data_0_in_valid = PENetwork_8_io_to_pes_0_in_valid; // @[pe.scala 264:34]
  assign PE_8_io_data_0_in_bits = PENetwork_8_io_to_pes_0_in_bits; // @[pe.scala 264:34]
  assign PE_9_clock = clock;
  assign PE_9_reset = reset;
  assign PE_9_io_data_2_sig_stat2trans = PENetwork_52_io_to_pes_9_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_9_io_data_1_in_valid = PENetwork_22_io_to_pes_9_in_valid; // @[pe.scala 264:34]
  assign PE_9_io_data_1_in_bits = PENetwork_22_io_to_pes_9_in_bits; // @[pe.scala 264:34]
  assign PE_9_io_data_0_in_valid = PENetwork_9_io_to_pes_0_in_valid; // @[pe.scala 264:34]
  assign PE_9_io_data_0_in_bits = PENetwork_9_io_to_pes_0_in_bits; // @[pe.scala 264:34]
  assign PE_10_clock = clock;
  assign PE_10_reset = reset;
  assign PE_10_io_data_2_sig_stat2trans = PENetwork_52_io_to_pes_10_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_10_io_data_1_in_valid = PENetwork_22_io_to_pes_10_in_valid; // @[pe.scala 264:34]
  assign PE_10_io_data_1_in_bits = PENetwork_22_io_to_pes_10_in_bits; // @[pe.scala 264:34]
  assign PE_10_io_data_0_in_valid = PENetwork_10_io_to_pes_0_in_valid; // @[pe.scala 264:34]
  assign PE_10_io_data_0_in_bits = PENetwork_10_io_to_pes_0_in_bits; // @[pe.scala 264:34]
  assign PE_11_clock = clock;
  assign PE_11_reset = reset;
  assign PE_11_io_data_2_sig_stat2trans = PENetwork_52_io_to_pes_11_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_11_io_data_1_in_valid = PENetwork_22_io_to_pes_11_in_valid; // @[pe.scala 264:34]
  assign PE_11_io_data_1_in_bits = PENetwork_22_io_to_pes_11_in_bits; // @[pe.scala 264:34]
  assign PE_11_io_data_0_in_valid = PENetwork_11_io_to_pes_0_in_valid; // @[pe.scala 264:34]
  assign PE_11_io_data_0_in_bits = PENetwork_11_io_to_pes_0_in_bits; // @[pe.scala 264:34]
  assign PE_12_clock = clock;
  assign PE_12_reset = reset;
  assign PE_12_io_data_2_sig_stat2trans = PENetwork_52_io_to_pes_12_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_12_io_data_1_in_valid = PENetwork_22_io_to_pes_12_in_valid; // @[pe.scala 264:34]
  assign PE_12_io_data_1_in_bits = PENetwork_22_io_to_pes_12_in_bits; // @[pe.scala 264:34]
  assign PE_12_io_data_0_in_valid = PENetwork_12_io_to_pes_0_in_valid; // @[pe.scala 264:34]
  assign PE_12_io_data_0_in_bits = PENetwork_12_io_to_pes_0_in_bits; // @[pe.scala 264:34]
  assign PE_13_clock = clock;
  assign PE_13_reset = reset;
  assign PE_13_io_data_2_sig_stat2trans = PENetwork_52_io_to_pes_13_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_13_io_data_1_in_valid = PENetwork_22_io_to_pes_13_in_valid; // @[pe.scala 264:34]
  assign PE_13_io_data_1_in_bits = PENetwork_22_io_to_pes_13_in_bits; // @[pe.scala 264:34]
  assign PE_13_io_data_0_in_valid = PENetwork_13_io_to_pes_0_in_valid; // @[pe.scala 264:34]
  assign PE_13_io_data_0_in_bits = PENetwork_13_io_to_pes_0_in_bits; // @[pe.scala 264:34]
  assign PE_14_clock = clock;
  assign PE_14_reset = reset;
  assign PE_14_io_data_2_sig_stat2trans = PENetwork_52_io_to_pes_14_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_14_io_data_1_in_valid = PENetwork_22_io_to_pes_14_in_valid; // @[pe.scala 264:34]
  assign PE_14_io_data_1_in_bits = PENetwork_22_io_to_pes_14_in_bits; // @[pe.scala 264:34]
  assign PE_14_io_data_0_in_valid = PENetwork_14_io_to_pes_0_in_valid; // @[pe.scala 264:34]
  assign PE_14_io_data_0_in_bits = PENetwork_14_io_to_pes_0_in_bits; // @[pe.scala 264:34]
  assign PE_15_clock = clock;
  assign PE_15_reset = reset;
  assign PE_15_io_data_2_sig_stat2trans = PENetwork_52_io_to_pes_15_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_15_io_data_1_in_valid = PENetwork_22_io_to_pes_15_in_valid; // @[pe.scala 264:34]
  assign PE_15_io_data_1_in_bits = PENetwork_22_io_to_pes_15_in_bits; // @[pe.scala 264:34]
  assign PE_15_io_data_0_in_valid = PENetwork_15_io_to_pes_0_in_valid; // @[pe.scala 264:34]
  assign PE_15_io_data_0_in_bits = PENetwork_15_io_to_pes_0_in_bits; // @[pe.scala 264:34]
  assign PE_16_clock = clock;
  assign PE_16_reset = reset;
  assign PE_16_io_data_2_sig_stat2trans = PENetwork_52_io_to_pes_16_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_16_io_data_1_in_valid = PENetwork_22_io_to_pes_16_in_valid; // @[pe.scala 264:34]
  assign PE_16_io_data_1_in_bits = PENetwork_22_io_to_pes_16_in_bits; // @[pe.scala 264:34]
  assign PE_16_io_data_0_in_valid = PENetwork_16_io_to_pes_0_in_valid; // @[pe.scala 264:34]
  assign PE_16_io_data_0_in_bits = PENetwork_16_io_to_pes_0_in_bits; // @[pe.scala 264:34]
  assign PE_17_clock = clock;
  assign PE_17_reset = reset;
  assign PE_17_io_data_2_sig_stat2trans = PENetwork_52_io_to_pes_17_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_17_io_data_1_in_valid = PENetwork_22_io_to_pes_17_in_valid; // @[pe.scala 264:34]
  assign PE_17_io_data_1_in_bits = PENetwork_22_io_to_pes_17_in_bits; // @[pe.scala 264:34]
  assign PE_17_io_data_0_in_valid = PENetwork_17_io_to_pes_0_in_valid; // @[pe.scala 264:34]
  assign PE_17_io_data_0_in_bits = PENetwork_17_io_to_pes_0_in_bits; // @[pe.scala 264:34]
  assign PE_18_clock = clock;
  assign PE_18_reset = reset;
  assign PE_18_io_data_2_sig_stat2trans = PENetwork_52_io_to_pes_18_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_18_io_data_1_in_valid = PENetwork_22_io_to_pes_18_in_valid; // @[pe.scala 264:34]
  assign PE_18_io_data_1_in_bits = PENetwork_22_io_to_pes_18_in_bits; // @[pe.scala 264:34]
  assign PE_18_io_data_0_in_valid = PENetwork_18_io_to_pes_0_in_valid; // @[pe.scala 264:34]
  assign PE_18_io_data_0_in_bits = PENetwork_18_io_to_pes_0_in_bits; // @[pe.scala 264:34]
  assign PE_19_clock = clock;
  assign PE_19_reset = reset;
  assign PE_19_io_data_2_sig_stat2trans = PENetwork_52_io_to_pes_19_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_19_io_data_1_in_valid = PENetwork_22_io_to_pes_19_in_valid; // @[pe.scala 264:34]
  assign PE_19_io_data_1_in_bits = PENetwork_22_io_to_pes_19_in_bits; // @[pe.scala 264:34]
  assign PE_19_io_data_0_in_valid = PENetwork_19_io_to_pes_0_in_valid; // @[pe.scala 264:34]
  assign PE_19_io_data_0_in_bits = PENetwork_19_io_to_pes_0_in_bits; // @[pe.scala 264:34]
  assign PE_20_clock = clock;
  assign PE_20_reset = reset;
  assign PE_20_io_data_2_sig_stat2trans = PENetwork_52_io_to_pes_20_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_20_io_data_1_in_valid = PENetwork_22_io_to_pes_20_in_valid; // @[pe.scala 264:34]
  assign PE_20_io_data_1_in_bits = PENetwork_22_io_to_pes_20_in_bits; // @[pe.scala 264:34]
  assign PE_20_io_data_0_in_valid = PENetwork_20_io_to_pes_0_in_valid; // @[pe.scala 264:34]
  assign PE_20_io_data_0_in_bits = PENetwork_20_io_to_pes_0_in_bits; // @[pe.scala 264:34]
  assign PE_21_clock = clock;
  assign PE_21_reset = reset;
  assign PE_21_io_data_2_sig_stat2trans = PENetwork_52_io_to_pes_21_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_21_io_data_1_in_valid = PENetwork_22_io_to_pes_21_in_valid; // @[pe.scala 264:34]
  assign PE_21_io_data_1_in_bits = PENetwork_22_io_to_pes_21_in_bits; // @[pe.scala 264:34]
  assign PE_21_io_data_0_in_valid = PENetwork_21_io_to_pes_0_in_valid; // @[pe.scala 264:34]
  assign PE_21_io_data_0_in_bits = PENetwork_21_io_to_pes_0_in_bits; // @[pe.scala 264:34]
  assign PE_22_clock = clock;
  assign PE_22_reset = reset;
  assign PE_22_io_data_2_sig_stat2trans = PENetwork_53_io_to_pes_0_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_22_io_data_1_in_valid = PENetwork_23_io_to_pes_0_in_valid; // @[pe.scala 264:34]
  assign PE_22_io_data_1_in_bits = PENetwork_23_io_to_pes_0_in_bits; // @[pe.scala 264:34]
  assign PE_22_io_data_0_in_valid = PENetwork_io_to_pes_1_in_valid; // @[pe.scala 264:34]
  assign PE_22_io_data_0_in_bits = PENetwork_io_to_pes_1_in_bits; // @[pe.scala 264:34]
  assign PE_23_clock = clock;
  assign PE_23_reset = reset;
  assign PE_23_io_data_2_sig_stat2trans = PENetwork_53_io_to_pes_1_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_23_io_data_1_in_valid = PENetwork_23_io_to_pes_1_in_valid; // @[pe.scala 264:34]
  assign PE_23_io_data_1_in_bits = PENetwork_23_io_to_pes_1_in_bits; // @[pe.scala 264:34]
  assign PE_23_io_data_0_in_valid = PENetwork_1_io_to_pes_1_in_valid; // @[pe.scala 264:34]
  assign PE_23_io_data_0_in_bits = PENetwork_1_io_to_pes_1_in_bits; // @[pe.scala 264:34]
  assign PE_24_clock = clock;
  assign PE_24_reset = reset;
  assign PE_24_io_data_2_sig_stat2trans = PENetwork_53_io_to_pes_2_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_24_io_data_1_in_valid = PENetwork_23_io_to_pes_2_in_valid; // @[pe.scala 264:34]
  assign PE_24_io_data_1_in_bits = PENetwork_23_io_to_pes_2_in_bits; // @[pe.scala 264:34]
  assign PE_24_io_data_0_in_valid = PENetwork_2_io_to_pes_1_in_valid; // @[pe.scala 264:34]
  assign PE_24_io_data_0_in_bits = PENetwork_2_io_to_pes_1_in_bits; // @[pe.scala 264:34]
  assign PE_25_clock = clock;
  assign PE_25_reset = reset;
  assign PE_25_io_data_2_sig_stat2trans = PENetwork_53_io_to_pes_3_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_25_io_data_1_in_valid = PENetwork_23_io_to_pes_3_in_valid; // @[pe.scala 264:34]
  assign PE_25_io_data_1_in_bits = PENetwork_23_io_to_pes_3_in_bits; // @[pe.scala 264:34]
  assign PE_25_io_data_0_in_valid = PENetwork_3_io_to_pes_1_in_valid; // @[pe.scala 264:34]
  assign PE_25_io_data_0_in_bits = PENetwork_3_io_to_pes_1_in_bits; // @[pe.scala 264:34]
  assign PE_26_clock = clock;
  assign PE_26_reset = reset;
  assign PE_26_io_data_2_sig_stat2trans = PENetwork_53_io_to_pes_4_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_26_io_data_1_in_valid = PENetwork_23_io_to_pes_4_in_valid; // @[pe.scala 264:34]
  assign PE_26_io_data_1_in_bits = PENetwork_23_io_to_pes_4_in_bits; // @[pe.scala 264:34]
  assign PE_26_io_data_0_in_valid = PENetwork_4_io_to_pes_1_in_valid; // @[pe.scala 264:34]
  assign PE_26_io_data_0_in_bits = PENetwork_4_io_to_pes_1_in_bits; // @[pe.scala 264:34]
  assign PE_27_clock = clock;
  assign PE_27_reset = reset;
  assign PE_27_io_data_2_sig_stat2trans = PENetwork_53_io_to_pes_5_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_27_io_data_1_in_valid = PENetwork_23_io_to_pes_5_in_valid; // @[pe.scala 264:34]
  assign PE_27_io_data_1_in_bits = PENetwork_23_io_to_pes_5_in_bits; // @[pe.scala 264:34]
  assign PE_27_io_data_0_in_valid = PENetwork_5_io_to_pes_1_in_valid; // @[pe.scala 264:34]
  assign PE_27_io_data_0_in_bits = PENetwork_5_io_to_pes_1_in_bits; // @[pe.scala 264:34]
  assign PE_28_clock = clock;
  assign PE_28_reset = reset;
  assign PE_28_io_data_2_sig_stat2trans = PENetwork_53_io_to_pes_6_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_28_io_data_1_in_valid = PENetwork_23_io_to_pes_6_in_valid; // @[pe.scala 264:34]
  assign PE_28_io_data_1_in_bits = PENetwork_23_io_to_pes_6_in_bits; // @[pe.scala 264:34]
  assign PE_28_io_data_0_in_valid = PENetwork_6_io_to_pes_1_in_valid; // @[pe.scala 264:34]
  assign PE_28_io_data_0_in_bits = PENetwork_6_io_to_pes_1_in_bits; // @[pe.scala 264:34]
  assign PE_29_clock = clock;
  assign PE_29_reset = reset;
  assign PE_29_io_data_2_sig_stat2trans = PENetwork_53_io_to_pes_7_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_29_io_data_1_in_valid = PENetwork_23_io_to_pes_7_in_valid; // @[pe.scala 264:34]
  assign PE_29_io_data_1_in_bits = PENetwork_23_io_to_pes_7_in_bits; // @[pe.scala 264:34]
  assign PE_29_io_data_0_in_valid = PENetwork_7_io_to_pes_1_in_valid; // @[pe.scala 264:34]
  assign PE_29_io_data_0_in_bits = PENetwork_7_io_to_pes_1_in_bits; // @[pe.scala 264:34]
  assign PE_30_clock = clock;
  assign PE_30_reset = reset;
  assign PE_30_io_data_2_sig_stat2trans = PENetwork_53_io_to_pes_8_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_30_io_data_1_in_valid = PENetwork_23_io_to_pes_8_in_valid; // @[pe.scala 264:34]
  assign PE_30_io_data_1_in_bits = PENetwork_23_io_to_pes_8_in_bits; // @[pe.scala 264:34]
  assign PE_30_io_data_0_in_valid = PENetwork_8_io_to_pes_1_in_valid; // @[pe.scala 264:34]
  assign PE_30_io_data_0_in_bits = PENetwork_8_io_to_pes_1_in_bits; // @[pe.scala 264:34]
  assign PE_31_clock = clock;
  assign PE_31_reset = reset;
  assign PE_31_io_data_2_sig_stat2trans = PENetwork_53_io_to_pes_9_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_31_io_data_1_in_valid = PENetwork_23_io_to_pes_9_in_valid; // @[pe.scala 264:34]
  assign PE_31_io_data_1_in_bits = PENetwork_23_io_to_pes_9_in_bits; // @[pe.scala 264:34]
  assign PE_31_io_data_0_in_valid = PENetwork_9_io_to_pes_1_in_valid; // @[pe.scala 264:34]
  assign PE_31_io_data_0_in_bits = PENetwork_9_io_to_pes_1_in_bits; // @[pe.scala 264:34]
  assign PE_32_clock = clock;
  assign PE_32_reset = reset;
  assign PE_32_io_data_2_sig_stat2trans = PENetwork_53_io_to_pes_10_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_32_io_data_1_in_valid = PENetwork_23_io_to_pes_10_in_valid; // @[pe.scala 264:34]
  assign PE_32_io_data_1_in_bits = PENetwork_23_io_to_pes_10_in_bits; // @[pe.scala 264:34]
  assign PE_32_io_data_0_in_valid = PENetwork_10_io_to_pes_1_in_valid; // @[pe.scala 264:34]
  assign PE_32_io_data_0_in_bits = PENetwork_10_io_to_pes_1_in_bits; // @[pe.scala 264:34]
  assign PE_33_clock = clock;
  assign PE_33_reset = reset;
  assign PE_33_io_data_2_sig_stat2trans = PENetwork_53_io_to_pes_11_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_33_io_data_1_in_valid = PENetwork_23_io_to_pes_11_in_valid; // @[pe.scala 264:34]
  assign PE_33_io_data_1_in_bits = PENetwork_23_io_to_pes_11_in_bits; // @[pe.scala 264:34]
  assign PE_33_io_data_0_in_valid = PENetwork_11_io_to_pes_1_in_valid; // @[pe.scala 264:34]
  assign PE_33_io_data_0_in_bits = PENetwork_11_io_to_pes_1_in_bits; // @[pe.scala 264:34]
  assign PE_34_clock = clock;
  assign PE_34_reset = reset;
  assign PE_34_io_data_2_sig_stat2trans = PENetwork_53_io_to_pes_12_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_34_io_data_1_in_valid = PENetwork_23_io_to_pes_12_in_valid; // @[pe.scala 264:34]
  assign PE_34_io_data_1_in_bits = PENetwork_23_io_to_pes_12_in_bits; // @[pe.scala 264:34]
  assign PE_34_io_data_0_in_valid = PENetwork_12_io_to_pes_1_in_valid; // @[pe.scala 264:34]
  assign PE_34_io_data_0_in_bits = PENetwork_12_io_to_pes_1_in_bits; // @[pe.scala 264:34]
  assign PE_35_clock = clock;
  assign PE_35_reset = reset;
  assign PE_35_io_data_2_sig_stat2trans = PENetwork_53_io_to_pes_13_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_35_io_data_1_in_valid = PENetwork_23_io_to_pes_13_in_valid; // @[pe.scala 264:34]
  assign PE_35_io_data_1_in_bits = PENetwork_23_io_to_pes_13_in_bits; // @[pe.scala 264:34]
  assign PE_35_io_data_0_in_valid = PENetwork_13_io_to_pes_1_in_valid; // @[pe.scala 264:34]
  assign PE_35_io_data_0_in_bits = PENetwork_13_io_to_pes_1_in_bits; // @[pe.scala 264:34]
  assign PE_36_clock = clock;
  assign PE_36_reset = reset;
  assign PE_36_io_data_2_sig_stat2trans = PENetwork_53_io_to_pes_14_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_36_io_data_1_in_valid = PENetwork_23_io_to_pes_14_in_valid; // @[pe.scala 264:34]
  assign PE_36_io_data_1_in_bits = PENetwork_23_io_to_pes_14_in_bits; // @[pe.scala 264:34]
  assign PE_36_io_data_0_in_valid = PENetwork_14_io_to_pes_1_in_valid; // @[pe.scala 264:34]
  assign PE_36_io_data_0_in_bits = PENetwork_14_io_to_pes_1_in_bits; // @[pe.scala 264:34]
  assign PE_37_clock = clock;
  assign PE_37_reset = reset;
  assign PE_37_io_data_2_sig_stat2trans = PENetwork_53_io_to_pes_15_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_37_io_data_1_in_valid = PENetwork_23_io_to_pes_15_in_valid; // @[pe.scala 264:34]
  assign PE_37_io_data_1_in_bits = PENetwork_23_io_to_pes_15_in_bits; // @[pe.scala 264:34]
  assign PE_37_io_data_0_in_valid = PENetwork_15_io_to_pes_1_in_valid; // @[pe.scala 264:34]
  assign PE_37_io_data_0_in_bits = PENetwork_15_io_to_pes_1_in_bits; // @[pe.scala 264:34]
  assign PE_38_clock = clock;
  assign PE_38_reset = reset;
  assign PE_38_io_data_2_sig_stat2trans = PENetwork_53_io_to_pes_16_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_38_io_data_1_in_valid = PENetwork_23_io_to_pes_16_in_valid; // @[pe.scala 264:34]
  assign PE_38_io_data_1_in_bits = PENetwork_23_io_to_pes_16_in_bits; // @[pe.scala 264:34]
  assign PE_38_io_data_0_in_valid = PENetwork_16_io_to_pes_1_in_valid; // @[pe.scala 264:34]
  assign PE_38_io_data_0_in_bits = PENetwork_16_io_to_pes_1_in_bits; // @[pe.scala 264:34]
  assign PE_39_clock = clock;
  assign PE_39_reset = reset;
  assign PE_39_io_data_2_sig_stat2trans = PENetwork_53_io_to_pes_17_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_39_io_data_1_in_valid = PENetwork_23_io_to_pes_17_in_valid; // @[pe.scala 264:34]
  assign PE_39_io_data_1_in_bits = PENetwork_23_io_to_pes_17_in_bits; // @[pe.scala 264:34]
  assign PE_39_io_data_0_in_valid = PENetwork_17_io_to_pes_1_in_valid; // @[pe.scala 264:34]
  assign PE_39_io_data_0_in_bits = PENetwork_17_io_to_pes_1_in_bits; // @[pe.scala 264:34]
  assign PE_40_clock = clock;
  assign PE_40_reset = reset;
  assign PE_40_io_data_2_sig_stat2trans = PENetwork_53_io_to_pes_18_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_40_io_data_1_in_valid = PENetwork_23_io_to_pes_18_in_valid; // @[pe.scala 264:34]
  assign PE_40_io_data_1_in_bits = PENetwork_23_io_to_pes_18_in_bits; // @[pe.scala 264:34]
  assign PE_40_io_data_0_in_valid = PENetwork_18_io_to_pes_1_in_valid; // @[pe.scala 264:34]
  assign PE_40_io_data_0_in_bits = PENetwork_18_io_to_pes_1_in_bits; // @[pe.scala 264:34]
  assign PE_41_clock = clock;
  assign PE_41_reset = reset;
  assign PE_41_io_data_2_sig_stat2trans = PENetwork_53_io_to_pes_19_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_41_io_data_1_in_valid = PENetwork_23_io_to_pes_19_in_valid; // @[pe.scala 264:34]
  assign PE_41_io_data_1_in_bits = PENetwork_23_io_to_pes_19_in_bits; // @[pe.scala 264:34]
  assign PE_41_io_data_0_in_valid = PENetwork_19_io_to_pes_1_in_valid; // @[pe.scala 264:34]
  assign PE_41_io_data_0_in_bits = PENetwork_19_io_to_pes_1_in_bits; // @[pe.scala 264:34]
  assign PE_42_clock = clock;
  assign PE_42_reset = reset;
  assign PE_42_io_data_2_sig_stat2trans = PENetwork_53_io_to_pes_20_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_42_io_data_1_in_valid = PENetwork_23_io_to_pes_20_in_valid; // @[pe.scala 264:34]
  assign PE_42_io_data_1_in_bits = PENetwork_23_io_to_pes_20_in_bits; // @[pe.scala 264:34]
  assign PE_42_io_data_0_in_valid = PENetwork_20_io_to_pes_1_in_valid; // @[pe.scala 264:34]
  assign PE_42_io_data_0_in_bits = PENetwork_20_io_to_pes_1_in_bits; // @[pe.scala 264:34]
  assign PE_43_clock = clock;
  assign PE_43_reset = reset;
  assign PE_43_io_data_2_sig_stat2trans = PENetwork_53_io_to_pes_21_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_43_io_data_1_in_valid = PENetwork_23_io_to_pes_21_in_valid; // @[pe.scala 264:34]
  assign PE_43_io_data_1_in_bits = PENetwork_23_io_to_pes_21_in_bits; // @[pe.scala 264:34]
  assign PE_43_io_data_0_in_valid = PENetwork_21_io_to_pes_1_in_valid; // @[pe.scala 264:34]
  assign PE_43_io_data_0_in_bits = PENetwork_21_io_to_pes_1_in_bits; // @[pe.scala 264:34]
  assign PE_44_clock = clock;
  assign PE_44_reset = reset;
  assign PE_44_io_data_2_sig_stat2trans = PENetwork_54_io_to_pes_0_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_44_io_data_1_in_valid = PENetwork_24_io_to_pes_0_in_valid; // @[pe.scala 264:34]
  assign PE_44_io_data_1_in_bits = PENetwork_24_io_to_pes_0_in_bits; // @[pe.scala 264:34]
  assign PE_44_io_data_0_in_valid = PENetwork_io_to_pes_2_in_valid; // @[pe.scala 264:34]
  assign PE_44_io_data_0_in_bits = PENetwork_io_to_pes_2_in_bits; // @[pe.scala 264:34]
  assign PE_45_clock = clock;
  assign PE_45_reset = reset;
  assign PE_45_io_data_2_sig_stat2trans = PENetwork_54_io_to_pes_1_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_45_io_data_1_in_valid = PENetwork_24_io_to_pes_1_in_valid; // @[pe.scala 264:34]
  assign PE_45_io_data_1_in_bits = PENetwork_24_io_to_pes_1_in_bits; // @[pe.scala 264:34]
  assign PE_45_io_data_0_in_valid = PENetwork_1_io_to_pes_2_in_valid; // @[pe.scala 264:34]
  assign PE_45_io_data_0_in_bits = PENetwork_1_io_to_pes_2_in_bits; // @[pe.scala 264:34]
  assign PE_46_clock = clock;
  assign PE_46_reset = reset;
  assign PE_46_io_data_2_sig_stat2trans = PENetwork_54_io_to_pes_2_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_46_io_data_1_in_valid = PENetwork_24_io_to_pes_2_in_valid; // @[pe.scala 264:34]
  assign PE_46_io_data_1_in_bits = PENetwork_24_io_to_pes_2_in_bits; // @[pe.scala 264:34]
  assign PE_46_io_data_0_in_valid = PENetwork_2_io_to_pes_2_in_valid; // @[pe.scala 264:34]
  assign PE_46_io_data_0_in_bits = PENetwork_2_io_to_pes_2_in_bits; // @[pe.scala 264:34]
  assign PE_47_clock = clock;
  assign PE_47_reset = reset;
  assign PE_47_io_data_2_sig_stat2trans = PENetwork_54_io_to_pes_3_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_47_io_data_1_in_valid = PENetwork_24_io_to_pes_3_in_valid; // @[pe.scala 264:34]
  assign PE_47_io_data_1_in_bits = PENetwork_24_io_to_pes_3_in_bits; // @[pe.scala 264:34]
  assign PE_47_io_data_0_in_valid = PENetwork_3_io_to_pes_2_in_valid; // @[pe.scala 264:34]
  assign PE_47_io_data_0_in_bits = PENetwork_3_io_to_pes_2_in_bits; // @[pe.scala 264:34]
  assign PE_48_clock = clock;
  assign PE_48_reset = reset;
  assign PE_48_io_data_2_sig_stat2trans = PENetwork_54_io_to_pes_4_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_48_io_data_1_in_valid = PENetwork_24_io_to_pes_4_in_valid; // @[pe.scala 264:34]
  assign PE_48_io_data_1_in_bits = PENetwork_24_io_to_pes_4_in_bits; // @[pe.scala 264:34]
  assign PE_48_io_data_0_in_valid = PENetwork_4_io_to_pes_2_in_valid; // @[pe.scala 264:34]
  assign PE_48_io_data_0_in_bits = PENetwork_4_io_to_pes_2_in_bits; // @[pe.scala 264:34]
  assign PE_49_clock = clock;
  assign PE_49_reset = reset;
  assign PE_49_io_data_2_sig_stat2trans = PENetwork_54_io_to_pes_5_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_49_io_data_1_in_valid = PENetwork_24_io_to_pes_5_in_valid; // @[pe.scala 264:34]
  assign PE_49_io_data_1_in_bits = PENetwork_24_io_to_pes_5_in_bits; // @[pe.scala 264:34]
  assign PE_49_io_data_0_in_valid = PENetwork_5_io_to_pes_2_in_valid; // @[pe.scala 264:34]
  assign PE_49_io_data_0_in_bits = PENetwork_5_io_to_pes_2_in_bits; // @[pe.scala 264:34]
  assign PE_50_clock = clock;
  assign PE_50_reset = reset;
  assign PE_50_io_data_2_sig_stat2trans = PENetwork_54_io_to_pes_6_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_50_io_data_1_in_valid = PENetwork_24_io_to_pes_6_in_valid; // @[pe.scala 264:34]
  assign PE_50_io_data_1_in_bits = PENetwork_24_io_to_pes_6_in_bits; // @[pe.scala 264:34]
  assign PE_50_io_data_0_in_valid = PENetwork_6_io_to_pes_2_in_valid; // @[pe.scala 264:34]
  assign PE_50_io_data_0_in_bits = PENetwork_6_io_to_pes_2_in_bits; // @[pe.scala 264:34]
  assign PE_51_clock = clock;
  assign PE_51_reset = reset;
  assign PE_51_io_data_2_sig_stat2trans = PENetwork_54_io_to_pes_7_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_51_io_data_1_in_valid = PENetwork_24_io_to_pes_7_in_valid; // @[pe.scala 264:34]
  assign PE_51_io_data_1_in_bits = PENetwork_24_io_to_pes_7_in_bits; // @[pe.scala 264:34]
  assign PE_51_io_data_0_in_valid = PENetwork_7_io_to_pes_2_in_valid; // @[pe.scala 264:34]
  assign PE_51_io_data_0_in_bits = PENetwork_7_io_to_pes_2_in_bits; // @[pe.scala 264:34]
  assign PE_52_clock = clock;
  assign PE_52_reset = reset;
  assign PE_52_io_data_2_sig_stat2trans = PENetwork_54_io_to_pes_8_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_52_io_data_1_in_valid = PENetwork_24_io_to_pes_8_in_valid; // @[pe.scala 264:34]
  assign PE_52_io_data_1_in_bits = PENetwork_24_io_to_pes_8_in_bits; // @[pe.scala 264:34]
  assign PE_52_io_data_0_in_valid = PENetwork_8_io_to_pes_2_in_valid; // @[pe.scala 264:34]
  assign PE_52_io_data_0_in_bits = PENetwork_8_io_to_pes_2_in_bits; // @[pe.scala 264:34]
  assign PE_53_clock = clock;
  assign PE_53_reset = reset;
  assign PE_53_io_data_2_sig_stat2trans = PENetwork_54_io_to_pes_9_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_53_io_data_1_in_valid = PENetwork_24_io_to_pes_9_in_valid; // @[pe.scala 264:34]
  assign PE_53_io_data_1_in_bits = PENetwork_24_io_to_pes_9_in_bits; // @[pe.scala 264:34]
  assign PE_53_io_data_0_in_valid = PENetwork_9_io_to_pes_2_in_valid; // @[pe.scala 264:34]
  assign PE_53_io_data_0_in_bits = PENetwork_9_io_to_pes_2_in_bits; // @[pe.scala 264:34]
  assign PE_54_clock = clock;
  assign PE_54_reset = reset;
  assign PE_54_io_data_2_sig_stat2trans = PENetwork_54_io_to_pes_10_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_54_io_data_1_in_valid = PENetwork_24_io_to_pes_10_in_valid; // @[pe.scala 264:34]
  assign PE_54_io_data_1_in_bits = PENetwork_24_io_to_pes_10_in_bits; // @[pe.scala 264:34]
  assign PE_54_io_data_0_in_valid = PENetwork_10_io_to_pes_2_in_valid; // @[pe.scala 264:34]
  assign PE_54_io_data_0_in_bits = PENetwork_10_io_to_pes_2_in_bits; // @[pe.scala 264:34]
  assign PE_55_clock = clock;
  assign PE_55_reset = reset;
  assign PE_55_io_data_2_sig_stat2trans = PENetwork_54_io_to_pes_11_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_55_io_data_1_in_valid = PENetwork_24_io_to_pes_11_in_valid; // @[pe.scala 264:34]
  assign PE_55_io_data_1_in_bits = PENetwork_24_io_to_pes_11_in_bits; // @[pe.scala 264:34]
  assign PE_55_io_data_0_in_valid = PENetwork_11_io_to_pes_2_in_valid; // @[pe.scala 264:34]
  assign PE_55_io_data_0_in_bits = PENetwork_11_io_to_pes_2_in_bits; // @[pe.scala 264:34]
  assign PE_56_clock = clock;
  assign PE_56_reset = reset;
  assign PE_56_io_data_2_sig_stat2trans = PENetwork_54_io_to_pes_12_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_56_io_data_1_in_valid = PENetwork_24_io_to_pes_12_in_valid; // @[pe.scala 264:34]
  assign PE_56_io_data_1_in_bits = PENetwork_24_io_to_pes_12_in_bits; // @[pe.scala 264:34]
  assign PE_56_io_data_0_in_valid = PENetwork_12_io_to_pes_2_in_valid; // @[pe.scala 264:34]
  assign PE_56_io_data_0_in_bits = PENetwork_12_io_to_pes_2_in_bits; // @[pe.scala 264:34]
  assign PE_57_clock = clock;
  assign PE_57_reset = reset;
  assign PE_57_io_data_2_sig_stat2trans = PENetwork_54_io_to_pes_13_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_57_io_data_1_in_valid = PENetwork_24_io_to_pes_13_in_valid; // @[pe.scala 264:34]
  assign PE_57_io_data_1_in_bits = PENetwork_24_io_to_pes_13_in_bits; // @[pe.scala 264:34]
  assign PE_57_io_data_0_in_valid = PENetwork_13_io_to_pes_2_in_valid; // @[pe.scala 264:34]
  assign PE_57_io_data_0_in_bits = PENetwork_13_io_to_pes_2_in_bits; // @[pe.scala 264:34]
  assign PE_58_clock = clock;
  assign PE_58_reset = reset;
  assign PE_58_io_data_2_sig_stat2trans = PENetwork_54_io_to_pes_14_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_58_io_data_1_in_valid = PENetwork_24_io_to_pes_14_in_valid; // @[pe.scala 264:34]
  assign PE_58_io_data_1_in_bits = PENetwork_24_io_to_pes_14_in_bits; // @[pe.scala 264:34]
  assign PE_58_io_data_0_in_valid = PENetwork_14_io_to_pes_2_in_valid; // @[pe.scala 264:34]
  assign PE_58_io_data_0_in_bits = PENetwork_14_io_to_pes_2_in_bits; // @[pe.scala 264:34]
  assign PE_59_clock = clock;
  assign PE_59_reset = reset;
  assign PE_59_io_data_2_sig_stat2trans = PENetwork_54_io_to_pes_15_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_59_io_data_1_in_valid = PENetwork_24_io_to_pes_15_in_valid; // @[pe.scala 264:34]
  assign PE_59_io_data_1_in_bits = PENetwork_24_io_to_pes_15_in_bits; // @[pe.scala 264:34]
  assign PE_59_io_data_0_in_valid = PENetwork_15_io_to_pes_2_in_valid; // @[pe.scala 264:34]
  assign PE_59_io_data_0_in_bits = PENetwork_15_io_to_pes_2_in_bits; // @[pe.scala 264:34]
  assign PE_60_clock = clock;
  assign PE_60_reset = reset;
  assign PE_60_io_data_2_sig_stat2trans = PENetwork_54_io_to_pes_16_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_60_io_data_1_in_valid = PENetwork_24_io_to_pes_16_in_valid; // @[pe.scala 264:34]
  assign PE_60_io_data_1_in_bits = PENetwork_24_io_to_pes_16_in_bits; // @[pe.scala 264:34]
  assign PE_60_io_data_0_in_valid = PENetwork_16_io_to_pes_2_in_valid; // @[pe.scala 264:34]
  assign PE_60_io_data_0_in_bits = PENetwork_16_io_to_pes_2_in_bits; // @[pe.scala 264:34]
  assign PE_61_clock = clock;
  assign PE_61_reset = reset;
  assign PE_61_io_data_2_sig_stat2trans = PENetwork_54_io_to_pes_17_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_61_io_data_1_in_valid = PENetwork_24_io_to_pes_17_in_valid; // @[pe.scala 264:34]
  assign PE_61_io_data_1_in_bits = PENetwork_24_io_to_pes_17_in_bits; // @[pe.scala 264:34]
  assign PE_61_io_data_0_in_valid = PENetwork_17_io_to_pes_2_in_valid; // @[pe.scala 264:34]
  assign PE_61_io_data_0_in_bits = PENetwork_17_io_to_pes_2_in_bits; // @[pe.scala 264:34]
  assign PE_62_clock = clock;
  assign PE_62_reset = reset;
  assign PE_62_io_data_2_sig_stat2trans = PENetwork_54_io_to_pes_18_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_62_io_data_1_in_valid = PENetwork_24_io_to_pes_18_in_valid; // @[pe.scala 264:34]
  assign PE_62_io_data_1_in_bits = PENetwork_24_io_to_pes_18_in_bits; // @[pe.scala 264:34]
  assign PE_62_io_data_0_in_valid = PENetwork_18_io_to_pes_2_in_valid; // @[pe.scala 264:34]
  assign PE_62_io_data_0_in_bits = PENetwork_18_io_to_pes_2_in_bits; // @[pe.scala 264:34]
  assign PE_63_clock = clock;
  assign PE_63_reset = reset;
  assign PE_63_io_data_2_sig_stat2trans = PENetwork_54_io_to_pes_19_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_63_io_data_1_in_valid = PENetwork_24_io_to_pes_19_in_valid; // @[pe.scala 264:34]
  assign PE_63_io_data_1_in_bits = PENetwork_24_io_to_pes_19_in_bits; // @[pe.scala 264:34]
  assign PE_63_io_data_0_in_valid = PENetwork_19_io_to_pes_2_in_valid; // @[pe.scala 264:34]
  assign PE_63_io_data_0_in_bits = PENetwork_19_io_to_pes_2_in_bits; // @[pe.scala 264:34]
  assign PE_64_clock = clock;
  assign PE_64_reset = reset;
  assign PE_64_io_data_2_sig_stat2trans = PENetwork_54_io_to_pes_20_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_64_io_data_1_in_valid = PENetwork_24_io_to_pes_20_in_valid; // @[pe.scala 264:34]
  assign PE_64_io_data_1_in_bits = PENetwork_24_io_to_pes_20_in_bits; // @[pe.scala 264:34]
  assign PE_64_io_data_0_in_valid = PENetwork_20_io_to_pes_2_in_valid; // @[pe.scala 264:34]
  assign PE_64_io_data_0_in_bits = PENetwork_20_io_to_pes_2_in_bits; // @[pe.scala 264:34]
  assign PE_65_clock = clock;
  assign PE_65_reset = reset;
  assign PE_65_io_data_2_sig_stat2trans = PENetwork_54_io_to_pes_21_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_65_io_data_1_in_valid = PENetwork_24_io_to_pes_21_in_valid; // @[pe.scala 264:34]
  assign PE_65_io_data_1_in_bits = PENetwork_24_io_to_pes_21_in_bits; // @[pe.scala 264:34]
  assign PE_65_io_data_0_in_valid = PENetwork_21_io_to_pes_2_in_valid; // @[pe.scala 264:34]
  assign PE_65_io_data_0_in_bits = PENetwork_21_io_to_pes_2_in_bits; // @[pe.scala 264:34]
  assign PE_66_clock = clock;
  assign PE_66_reset = reset;
  assign PE_66_io_data_2_sig_stat2trans = PENetwork_55_io_to_pes_0_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_66_io_data_1_in_valid = PENetwork_25_io_to_pes_0_in_valid; // @[pe.scala 264:34]
  assign PE_66_io_data_1_in_bits = PENetwork_25_io_to_pes_0_in_bits; // @[pe.scala 264:34]
  assign PE_66_io_data_0_in_valid = PENetwork_io_to_pes_3_in_valid; // @[pe.scala 264:34]
  assign PE_66_io_data_0_in_bits = PENetwork_io_to_pes_3_in_bits; // @[pe.scala 264:34]
  assign PE_67_clock = clock;
  assign PE_67_reset = reset;
  assign PE_67_io_data_2_sig_stat2trans = PENetwork_55_io_to_pes_1_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_67_io_data_1_in_valid = PENetwork_25_io_to_pes_1_in_valid; // @[pe.scala 264:34]
  assign PE_67_io_data_1_in_bits = PENetwork_25_io_to_pes_1_in_bits; // @[pe.scala 264:34]
  assign PE_67_io_data_0_in_valid = PENetwork_1_io_to_pes_3_in_valid; // @[pe.scala 264:34]
  assign PE_67_io_data_0_in_bits = PENetwork_1_io_to_pes_3_in_bits; // @[pe.scala 264:34]
  assign PE_68_clock = clock;
  assign PE_68_reset = reset;
  assign PE_68_io_data_2_sig_stat2trans = PENetwork_55_io_to_pes_2_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_68_io_data_1_in_valid = PENetwork_25_io_to_pes_2_in_valid; // @[pe.scala 264:34]
  assign PE_68_io_data_1_in_bits = PENetwork_25_io_to_pes_2_in_bits; // @[pe.scala 264:34]
  assign PE_68_io_data_0_in_valid = PENetwork_2_io_to_pes_3_in_valid; // @[pe.scala 264:34]
  assign PE_68_io_data_0_in_bits = PENetwork_2_io_to_pes_3_in_bits; // @[pe.scala 264:34]
  assign PE_69_clock = clock;
  assign PE_69_reset = reset;
  assign PE_69_io_data_2_sig_stat2trans = PENetwork_55_io_to_pes_3_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_69_io_data_1_in_valid = PENetwork_25_io_to_pes_3_in_valid; // @[pe.scala 264:34]
  assign PE_69_io_data_1_in_bits = PENetwork_25_io_to_pes_3_in_bits; // @[pe.scala 264:34]
  assign PE_69_io_data_0_in_valid = PENetwork_3_io_to_pes_3_in_valid; // @[pe.scala 264:34]
  assign PE_69_io_data_0_in_bits = PENetwork_3_io_to_pes_3_in_bits; // @[pe.scala 264:34]
  assign PE_70_clock = clock;
  assign PE_70_reset = reset;
  assign PE_70_io_data_2_sig_stat2trans = PENetwork_55_io_to_pes_4_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_70_io_data_1_in_valid = PENetwork_25_io_to_pes_4_in_valid; // @[pe.scala 264:34]
  assign PE_70_io_data_1_in_bits = PENetwork_25_io_to_pes_4_in_bits; // @[pe.scala 264:34]
  assign PE_70_io_data_0_in_valid = PENetwork_4_io_to_pes_3_in_valid; // @[pe.scala 264:34]
  assign PE_70_io_data_0_in_bits = PENetwork_4_io_to_pes_3_in_bits; // @[pe.scala 264:34]
  assign PE_71_clock = clock;
  assign PE_71_reset = reset;
  assign PE_71_io_data_2_sig_stat2trans = PENetwork_55_io_to_pes_5_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_71_io_data_1_in_valid = PENetwork_25_io_to_pes_5_in_valid; // @[pe.scala 264:34]
  assign PE_71_io_data_1_in_bits = PENetwork_25_io_to_pes_5_in_bits; // @[pe.scala 264:34]
  assign PE_71_io_data_0_in_valid = PENetwork_5_io_to_pes_3_in_valid; // @[pe.scala 264:34]
  assign PE_71_io_data_0_in_bits = PENetwork_5_io_to_pes_3_in_bits; // @[pe.scala 264:34]
  assign PE_72_clock = clock;
  assign PE_72_reset = reset;
  assign PE_72_io_data_2_sig_stat2trans = PENetwork_55_io_to_pes_6_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_72_io_data_1_in_valid = PENetwork_25_io_to_pes_6_in_valid; // @[pe.scala 264:34]
  assign PE_72_io_data_1_in_bits = PENetwork_25_io_to_pes_6_in_bits; // @[pe.scala 264:34]
  assign PE_72_io_data_0_in_valid = PENetwork_6_io_to_pes_3_in_valid; // @[pe.scala 264:34]
  assign PE_72_io_data_0_in_bits = PENetwork_6_io_to_pes_3_in_bits; // @[pe.scala 264:34]
  assign PE_73_clock = clock;
  assign PE_73_reset = reset;
  assign PE_73_io_data_2_sig_stat2trans = PENetwork_55_io_to_pes_7_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_73_io_data_1_in_valid = PENetwork_25_io_to_pes_7_in_valid; // @[pe.scala 264:34]
  assign PE_73_io_data_1_in_bits = PENetwork_25_io_to_pes_7_in_bits; // @[pe.scala 264:34]
  assign PE_73_io_data_0_in_valid = PENetwork_7_io_to_pes_3_in_valid; // @[pe.scala 264:34]
  assign PE_73_io_data_0_in_bits = PENetwork_7_io_to_pes_3_in_bits; // @[pe.scala 264:34]
  assign PE_74_clock = clock;
  assign PE_74_reset = reset;
  assign PE_74_io_data_2_sig_stat2trans = PENetwork_55_io_to_pes_8_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_74_io_data_1_in_valid = PENetwork_25_io_to_pes_8_in_valid; // @[pe.scala 264:34]
  assign PE_74_io_data_1_in_bits = PENetwork_25_io_to_pes_8_in_bits; // @[pe.scala 264:34]
  assign PE_74_io_data_0_in_valid = PENetwork_8_io_to_pes_3_in_valid; // @[pe.scala 264:34]
  assign PE_74_io_data_0_in_bits = PENetwork_8_io_to_pes_3_in_bits; // @[pe.scala 264:34]
  assign PE_75_clock = clock;
  assign PE_75_reset = reset;
  assign PE_75_io_data_2_sig_stat2trans = PENetwork_55_io_to_pes_9_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_75_io_data_1_in_valid = PENetwork_25_io_to_pes_9_in_valid; // @[pe.scala 264:34]
  assign PE_75_io_data_1_in_bits = PENetwork_25_io_to_pes_9_in_bits; // @[pe.scala 264:34]
  assign PE_75_io_data_0_in_valid = PENetwork_9_io_to_pes_3_in_valid; // @[pe.scala 264:34]
  assign PE_75_io_data_0_in_bits = PENetwork_9_io_to_pes_3_in_bits; // @[pe.scala 264:34]
  assign PE_76_clock = clock;
  assign PE_76_reset = reset;
  assign PE_76_io_data_2_sig_stat2trans = PENetwork_55_io_to_pes_10_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_76_io_data_1_in_valid = PENetwork_25_io_to_pes_10_in_valid; // @[pe.scala 264:34]
  assign PE_76_io_data_1_in_bits = PENetwork_25_io_to_pes_10_in_bits; // @[pe.scala 264:34]
  assign PE_76_io_data_0_in_valid = PENetwork_10_io_to_pes_3_in_valid; // @[pe.scala 264:34]
  assign PE_76_io_data_0_in_bits = PENetwork_10_io_to_pes_3_in_bits; // @[pe.scala 264:34]
  assign PE_77_clock = clock;
  assign PE_77_reset = reset;
  assign PE_77_io_data_2_sig_stat2trans = PENetwork_55_io_to_pes_11_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_77_io_data_1_in_valid = PENetwork_25_io_to_pes_11_in_valid; // @[pe.scala 264:34]
  assign PE_77_io_data_1_in_bits = PENetwork_25_io_to_pes_11_in_bits; // @[pe.scala 264:34]
  assign PE_77_io_data_0_in_valid = PENetwork_11_io_to_pes_3_in_valid; // @[pe.scala 264:34]
  assign PE_77_io_data_0_in_bits = PENetwork_11_io_to_pes_3_in_bits; // @[pe.scala 264:34]
  assign PE_78_clock = clock;
  assign PE_78_reset = reset;
  assign PE_78_io_data_2_sig_stat2trans = PENetwork_55_io_to_pes_12_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_78_io_data_1_in_valid = PENetwork_25_io_to_pes_12_in_valid; // @[pe.scala 264:34]
  assign PE_78_io_data_1_in_bits = PENetwork_25_io_to_pes_12_in_bits; // @[pe.scala 264:34]
  assign PE_78_io_data_0_in_valid = PENetwork_12_io_to_pes_3_in_valid; // @[pe.scala 264:34]
  assign PE_78_io_data_0_in_bits = PENetwork_12_io_to_pes_3_in_bits; // @[pe.scala 264:34]
  assign PE_79_clock = clock;
  assign PE_79_reset = reset;
  assign PE_79_io_data_2_sig_stat2trans = PENetwork_55_io_to_pes_13_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_79_io_data_1_in_valid = PENetwork_25_io_to_pes_13_in_valid; // @[pe.scala 264:34]
  assign PE_79_io_data_1_in_bits = PENetwork_25_io_to_pes_13_in_bits; // @[pe.scala 264:34]
  assign PE_79_io_data_0_in_valid = PENetwork_13_io_to_pes_3_in_valid; // @[pe.scala 264:34]
  assign PE_79_io_data_0_in_bits = PENetwork_13_io_to_pes_3_in_bits; // @[pe.scala 264:34]
  assign PE_80_clock = clock;
  assign PE_80_reset = reset;
  assign PE_80_io_data_2_sig_stat2trans = PENetwork_55_io_to_pes_14_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_80_io_data_1_in_valid = PENetwork_25_io_to_pes_14_in_valid; // @[pe.scala 264:34]
  assign PE_80_io_data_1_in_bits = PENetwork_25_io_to_pes_14_in_bits; // @[pe.scala 264:34]
  assign PE_80_io_data_0_in_valid = PENetwork_14_io_to_pes_3_in_valid; // @[pe.scala 264:34]
  assign PE_80_io_data_0_in_bits = PENetwork_14_io_to_pes_3_in_bits; // @[pe.scala 264:34]
  assign PE_81_clock = clock;
  assign PE_81_reset = reset;
  assign PE_81_io_data_2_sig_stat2trans = PENetwork_55_io_to_pes_15_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_81_io_data_1_in_valid = PENetwork_25_io_to_pes_15_in_valid; // @[pe.scala 264:34]
  assign PE_81_io_data_1_in_bits = PENetwork_25_io_to_pes_15_in_bits; // @[pe.scala 264:34]
  assign PE_81_io_data_0_in_valid = PENetwork_15_io_to_pes_3_in_valid; // @[pe.scala 264:34]
  assign PE_81_io_data_0_in_bits = PENetwork_15_io_to_pes_3_in_bits; // @[pe.scala 264:34]
  assign PE_82_clock = clock;
  assign PE_82_reset = reset;
  assign PE_82_io_data_2_sig_stat2trans = PENetwork_55_io_to_pes_16_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_82_io_data_1_in_valid = PENetwork_25_io_to_pes_16_in_valid; // @[pe.scala 264:34]
  assign PE_82_io_data_1_in_bits = PENetwork_25_io_to_pes_16_in_bits; // @[pe.scala 264:34]
  assign PE_82_io_data_0_in_valid = PENetwork_16_io_to_pes_3_in_valid; // @[pe.scala 264:34]
  assign PE_82_io_data_0_in_bits = PENetwork_16_io_to_pes_3_in_bits; // @[pe.scala 264:34]
  assign PE_83_clock = clock;
  assign PE_83_reset = reset;
  assign PE_83_io_data_2_sig_stat2trans = PENetwork_55_io_to_pes_17_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_83_io_data_1_in_valid = PENetwork_25_io_to_pes_17_in_valid; // @[pe.scala 264:34]
  assign PE_83_io_data_1_in_bits = PENetwork_25_io_to_pes_17_in_bits; // @[pe.scala 264:34]
  assign PE_83_io_data_0_in_valid = PENetwork_17_io_to_pes_3_in_valid; // @[pe.scala 264:34]
  assign PE_83_io_data_0_in_bits = PENetwork_17_io_to_pes_3_in_bits; // @[pe.scala 264:34]
  assign PE_84_clock = clock;
  assign PE_84_reset = reset;
  assign PE_84_io_data_2_sig_stat2trans = PENetwork_55_io_to_pes_18_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_84_io_data_1_in_valid = PENetwork_25_io_to_pes_18_in_valid; // @[pe.scala 264:34]
  assign PE_84_io_data_1_in_bits = PENetwork_25_io_to_pes_18_in_bits; // @[pe.scala 264:34]
  assign PE_84_io_data_0_in_valid = PENetwork_18_io_to_pes_3_in_valid; // @[pe.scala 264:34]
  assign PE_84_io_data_0_in_bits = PENetwork_18_io_to_pes_3_in_bits; // @[pe.scala 264:34]
  assign PE_85_clock = clock;
  assign PE_85_reset = reset;
  assign PE_85_io_data_2_sig_stat2trans = PENetwork_55_io_to_pes_19_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_85_io_data_1_in_valid = PENetwork_25_io_to_pes_19_in_valid; // @[pe.scala 264:34]
  assign PE_85_io_data_1_in_bits = PENetwork_25_io_to_pes_19_in_bits; // @[pe.scala 264:34]
  assign PE_85_io_data_0_in_valid = PENetwork_19_io_to_pes_3_in_valid; // @[pe.scala 264:34]
  assign PE_85_io_data_0_in_bits = PENetwork_19_io_to_pes_3_in_bits; // @[pe.scala 264:34]
  assign PE_86_clock = clock;
  assign PE_86_reset = reset;
  assign PE_86_io_data_2_sig_stat2trans = PENetwork_55_io_to_pes_20_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_86_io_data_1_in_valid = PENetwork_25_io_to_pes_20_in_valid; // @[pe.scala 264:34]
  assign PE_86_io_data_1_in_bits = PENetwork_25_io_to_pes_20_in_bits; // @[pe.scala 264:34]
  assign PE_86_io_data_0_in_valid = PENetwork_20_io_to_pes_3_in_valid; // @[pe.scala 264:34]
  assign PE_86_io_data_0_in_bits = PENetwork_20_io_to_pes_3_in_bits; // @[pe.scala 264:34]
  assign PE_87_clock = clock;
  assign PE_87_reset = reset;
  assign PE_87_io_data_2_sig_stat2trans = PENetwork_55_io_to_pes_21_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_87_io_data_1_in_valid = PENetwork_25_io_to_pes_21_in_valid; // @[pe.scala 264:34]
  assign PE_87_io_data_1_in_bits = PENetwork_25_io_to_pes_21_in_bits; // @[pe.scala 264:34]
  assign PE_87_io_data_0_in_valid = PENetwork_21_io_to_pes_3_in_valid; // @[pe.scala 264:34]
  assign PE_87_io_data_0_in_bits = PENetwork_21_io_to_pes_3_in_bits; // @[pe.scala 264:34]
  assign PE_88_clock = clock;
  assign PE_88_reset = reset;
  assign PE_88_io_data_2_sig_stat2trans = PENetwork_56_io_to_pes_0_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_88_io_data_1_in_valid = PENetwork_26_io_to_pes_0_in_valid; // @[pe.scala 264:34]
  assign PE_88_io_data_1_in_bits = PENetwork_26_io_to_pes_0_in_bits; // @[pe.scala 264:34]
  assign PE_88_io_data_0_in_valid = PENetwork_io_to_pes_4_in_valid; // @[pe.scala 264:34]
  assign PE_88_io_data_0_in_bits = PENetwork_io_to_pes_4_in_bits; // @[pe.scala 264:34]
  assign PE_89_clock = clock;
  assign PE_89_reset = reset;
  assign PE_89_io_data_2_sig_stat2trans = PENetwork_56_io_to_pes_1_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_89_io_data_1_in_valid = PENetwork_26_io_to_pes_1_in_valid; // @[pe.scala 264:34]
  assign PE_89_io_data_1_in_bits = PENetwork_26_io_to_pes_1_in_bits; // @[pe.scala 264:34]
  assign PE_89_io_data_0_in_valid = PENetwork_1_io_to_pes_4_in_valid; // @[pe.scala 264:34]
  assign PE_89_io_data_0_in_bits = PENetwork_1_io_to_pes_4_in_bits; // @[pe.scala 264:34]
  assign PE_90_clock = clock;
  assign PE_90_reset = reset;
  assign PE_90_io_data_2_sig_stat2trans = PENetwork_56_io_to_pes_2_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_90_io_data_1_in_valid = PENetwork_26_io_to_pes_2_in_valid; // @[pe.scala 264:34]
  assign PE_90_io_data_1_in_bits = PENetwork_26_io_to_pes_2_in_bits; // @[pe.scala 264:34]
  assign PE_90_io_data_0_in_valid = PENetwork_2_io_to_pes_4_in_valid; // @[pe.scala 264:34]
  assign PE_90_io_data_0_in_bits = PENetwork_2_io_to_pes_4_in_bits; // @[pe.scala 264:34]
  assign PE_91_clock = clock;
  assign PE_91_reset = reset;
  assign PE_91_io_data_2_sig_stat2trans = PENetwork_56_io_to_pes_3_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_91_io_data_1_in_valid = PENetwork_26_io_to_pes_3_in_valid; // @[pe.scala 264:34]
  assign PE_91_io_data_1_in_bits = PENetwork_26_io_to_pes_3_in_bits; // @[pe.scala 264:34]
  assign PE_91_io_data_0_in_valid = PENetwork_3_io_to_pes_4_in_valid; // @[pe.scala 264:34]
  assign PE_91_io_data_0_in_bits = PENetwork_3_io_to_pes_4_in_bits; // @[pe.scala 264:34]
  assign PE_92_clock = clock;
  assign PE_92_reset = reset;
  assign PE_92_io_data_2_sig_stat2trans = PENetwork_56_io_to_pes_4_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_92_io_data_1_in_valid = PENetwork_26_io_to_pes_4_in_valid; // @[pe.scala 264:34]
  assign PE_92_io_data_1_in_bits = PENetwork_26_io_to_pes_4_in_bits; // @[pe.scala 264:34]
  assign PE_92_io_data_0_in_valid = PENetwork_4_io_to_pes_4_in_valid; // @[pe.scala 264:34]
  assign PE_92_io_data_0_in_bits = PENetwork_4_io_to_pes_4_in_bits; // @[pe.scala 264:34]
  assign PE_93_clock = clock;
  assign PE_93_reset = reset;
  assign PE_93_io_data_2_sig_stat2trans = PENetwork_56_io_to_pes_5_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_93_io_data_1_in_valid = PENetwork_26_io_to_pes_5_in_valid; // @[pe.scala 264:34]
  assign PE_93_io_data_1_in_bits = PENetwork_26_io_to_pes_5_in_bits; // @[pe.scala 264:34]
  assign PE_93_io_data_0_in_valid = PENetwork_5_io_to_pes_4_in_valid; // @[pe.scala 264:34]
  assign PE_93_io_data_0_in_bits = PENetwork_5_io_to_pes_4_in_bits; // @[pe.scala 264:34]
  assign PE_94_clock = clock;
  assign PE_94_reset = reset;
  assign PE_94_io_data_2_sig_stat2trans = PENetwork_56_io_to_pes_6_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_94_io_data_1_in_valid = PENetwork_26_io_to_pes_6_in_valid; // @[pe.scala 264:34]
  assign PE_94_io_data_1_in_bits = PENetwork_26_io_to_pes_6_in_bits; // @[pe.scala 264:34]
  assign PE_94_io_data_0_in_valid = PENetwork_6_io_to_pes_4_in_valid; // @[pe.scala 264:34]
  assign PE_94_io_data_0_in_bits = PENetwork_6_io_to_pes_4_in_bits; // @[pe.scala 264:34]
  assign PE_95_clock = clock;
  assign PE_95_reset = reset;
  assign PE_95_io_data_2_sig_stat2trans = PENetwork_56_io_to_pes_7_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_95_io_data_1_in_valid = PENetwork_26_io_to_pes_7_in_valid; // @[pe.scala 264:34]
  assign PE_95_io_data_1_in_bits = PENetwork_26_io_to_pes_7_in_bits; // @[pe.scala 264:34]
  assign PE_95_io_data_0_in_valid = PENetwork_7_io_to_pes_4_in_valid; // @[pe.scala 264:34]
  assign PE_95_io_data_0_in_bits = PENetwork_7_io_to_pes_4_in_bits; // @[pe.scala 264:34]
  assign PE_96_clock = clock;
  assign PE_96_reset = reset;
  assign PE_96_io_data_2_sig_stat2trans = PENetwork_56_io_to_pes_8_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_96_io_data_1_in_valid = PENetwork_26_io_to_pes_8_in_valid; // @[pe.scala 264:34]
  assign PE_96_io_data_1_in_bits = PENetwork_26_io_to_pes_8_in_bits; // @[pe.scala 264:34]
  assign PE_96_io_data_0_in_valid = PENetwork_8_io_to_pes_4_in_valid; // @[pe.scala 264:34]
  assign PE_96_io_data_0_in_bits = PENetwork_8_io_to_pes_4_in_bits; // @[pe.scala 264:34]
  assign PE_97_clock = clock;
  assign PE_97_reset = reset;
  assign PE_97_io_data_2_sig_stat2trans = PENetwork_56_io_to_pes_9_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_97_io_data_1_in_valid = PENetwork_26_io_to_pes_9_in_valid; // @[pe.scala 264:34]
  assign PE_97_io_data_1_in_bits = PENetwork_26_io_to_pes_9_in_bits; // @[pe.scala 264:34]
  assign PE_97_io_data_0_in_valid = PENetwork_9_io_to_pes_4_in_valid; // @[pe.scala 264:34]
  assign PE_97_io_data_0_in_bits = PENetwork_9_io_to_pes_4_in_bits; // @[pe.scala 264:34]
  assign PE_98_clock = clock;
  assign PE_98_reset = reset;
  assign PE_98_io_data_2_sig_stat2trans = PENetwork_56_io_to_pes_10_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_98_io_data_1_in_valid = PENetwork_26_io_to_pes_10_in_valid; // @[pe.scala 264:34]
  assign PE_98_io_data_1_in_bits = PENetwork_26_io_to_pes_10_in_bits; // @[pe.scala 264:34]
  assign PE_98_io_data_0_in_valid = PENetwork_10_io_to_pes_4_in_valid; // @[pe.scala 264:34]
  assign PE_98_io_data_0_in_bits = PENetwork_10_io_to_pes_4_in_bits; // @[pe.scala 264:34]
  assign PE_99_clock = clock;
  assign PE_99_reset = reset;
  assign PE_99_io_data_2_sig_stat2trans = PENetwork_56_io_to_pes_11_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_99_io_data_1_in_valid = PENetwork_26_io_to_pes_11_in_valid; // @[pe.scala 264:34]
  assign PE_99_io_data_1_in_bits = PENetwork_26_io_to_pes_11_in_bits; // @[pe.scala 264:34]
  assign PE_99_io_data_0_in_valid = PENetwork_11_io_to_pes_4_in_valid; // @[pe.scala 264:34]
  assign PE_99_io_data_0_in_bits = PENetwork_11_io_to_pes_4_in_bits; // @[pe.scala 264:34]
  assign PE_100_clock = clock;
  assign PE_100_reset = reset;
  assign PE_100_io_data_2_sig_stat2trans = PENetwork_56_io_to_pes_12_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_100_io_data_1_in_valid = PENetwork_26_io_to_pes_12_in_valid; // @[pe.scala 264:34]
  assign PE_100_io_data_1_in_bits = PENetwork_26_io_to_pes_12_in_bits; // @[pe.scala 264:34]
  assign PE_100_io_data_0_in_valid = PENetwork_12_io_to_pes_4_in_valid; // @[pe.scala 264:34]
  assign PE_100_io_data_0_in_bits = PENetwork_12_io_to_pes_4_in_bits; // @[pe.scala 264:34]
  assign PE_101_clock = clock;
  assign PE_101_reset = reset;
  assign PE_101_io_data_2_sig_stat2trans = PENetwork_56_io_to_pes_13_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_101_io_data_1_in_valid = PENetwork_26_io_to_pes_13_in_valid; // @[pe.scala 264:34]
  assign PE_101_io_data_1_in_bits = PENetwork_26_io_to_pes_13_in_bits; // @[pe.scala 264:34]
  assign PE_101_io_data_0_in_valid = PENetwork_13_io_to_pes_4_in_valid; // @[pe.scala 264:34]
  assign PE_101_io_data_0_in_bits = PENetwork_13_io_to_pes_4_in_bits; // @[pe.scala 264:34]
  assign PE_102_clock = clock;
  assign PE_102_reset = reset;
  assign PE_102_io_data_2_sig_stat2trans = PENetwork_56_io_to_pes_14_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_102_io_data_1_in_valid = PENetwork_26_io_to_pes_14_in_valid; // @[pe.scala 264:34]
  assign PE_102_io_data_1_in_bits = PENetwork_26_io_to_pes_14_in_bits; // @[pe.scala 264:34]
  assign PE_102_io_data_0_in_valid = PENetwork_14_io_to_pes_4_in_valid; // @[pe.scala 264:34]
  assign PE_102_io_data_0_in_bits = PENetwork_14_io_to_pes_4_in_bits; // @[pe.scala 264:34]
  assign PE_103_clock = clock;
  assign PE_103_reset = reset;
  assign PE_103_io_data_2_sig_stat2trans = PENetwork_56_io_to_pes_15_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_103_io_data_1_in_valid = PENetwork_26_io_to_pes_15_in_valid; // @[pe.scala 264:34]
  assign PE_103_io_data_1_in_bits = PENetwork_26_io_to_pes_15_in_bits; // @[pe.scala 264:34]
  assign PE_103_io_data_0_in_valid = PENetwork_15_io_to_pes_4_in_valid; // @[pe.scala 264:34]
  assign PE_103_io_data_0_in_bits = PENetwork_15_io_to_pes_4_in_bits; // @[pe.scala 264:34]
  assign PE_104_clock = clock;
  assign PE_104_reset = reset;
  assign PE_104_io_data_2_sig_stat2trans = PENetwork_56_io_to_pes_16_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_104_io_data_1_in_valid = PENetwork_26_io_to_pes_16_in_valid; // @[pe.scala 264:34]
  assign PE_104_io_data_1_in_bits = PENetwork_26_io_to_pes_16_in_bits; // @[pe.scala 264:34]
  assign PE_104_io_data_0_in_valid = PENetwork_16_io_to_pes_4_in_valid; // @[pe.scala 264:34]
  assign PE_104_io_data_0_in_bits = PENetwork_16_io_to_pes_4_in_bits; // @[pe.scala 264:34]
  assign PE_105_clock = clock;
  assign PE_105_reset = reset;
  assign PE_105_io_data_2_sig_stat2trans = PENetwork_56_io_to_pes_17_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_105_io_data_1_in_valid = PENetwork_26_io_to_pes_17_in_valid; // @[pe.scala 264:34]
  assign PE_105_io_data_1_in_bits = PENetwork_26_io_to_pes_17_in_bits; // @[pe.scala 264:34]
  assign PE_105_io_data_0_in_valid = PENetwork_17_io_to_pes_4_in_valid; // @[pe.scala 264:34]
  assign PE_105_io_data_0_in_bits = PENetwork_17_io_to_pes_4_in_bits; // @[pe.scala 264:34]
  assign PE_106_clock = clock;
  assign PE_106_reset = reset;
  assign PE_106_io_data_2_sig_stat2trans = PENetwork_56_io_to_pes_18_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_106_io_data_1_in_valid = PENetwork_26_io_to_pes_18_in_valid; // @[pe.scala 264:34]
  assign PE_106_io_data_1_in_bits = PENetwork_26_io_to_pes_18_in_bits; // @[pe.scala 264:34]
  assign PE_106_io_data_0_in_valid = PENetwork_18_io_to_pes_4_in_valid; // @[pe.scala 264:34]
  assign PE_106_io_data_0_in_bits = PENetwork_18_io_to_pes_4_in_bits; // @[pe.scala 264:34]
  assign PE_107_clock = clock;
  assign PE_107_reset = reset;
  assign PE_107_io_data_2_sig_stat2trans = PENetwork_56_io_to_pes_19_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_107_io_data_1_in_valid = PENetwork_26_io_to_pes_19_in_valid; // @[pe.scala 264:34]
  assign PE_107_io_data_1_in_bits = PENetwork_26_io_to_pes_19_in_bits; // @[pe.scala 264:34]
  assign PE_107_io_data_0_in_valid = PENetwork_19_io_to_pes_4_in_valid; // @[pe.scala 264:34]
  assign PE_107_io_data_0_in_bits = PENetwork_19_io_to_pes_4_in_bits; // @[pe.scala 264:34]
  assign PE_108_clock = clock;
  assign PE_108_reset = reset;
  assign PE_108_io_data_2_sig_stat2trans = PENetwork_56_io_to_pes_20_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_108_io_data_1_in_valid = PENetwork_26_io_to_pes_20_in_valid; // @[pe.scala 264:34]
  assign PE_108_io_data_1_in_bits = PENetwork_26_io_to_pes_20_in_bits; // @[pe.scala 264:34]
  assign PE_108_io_data_0_in_valid = PENetwork_20_io_to_pes_4_in_valid; // @[pe.scala 264:34]
  assign PE_108_io_data_0_in_bits = PENetwork_20_io_to_pes_4_in_bits; // @[pe.scala 264:34]
  assign PE_109_clock = clock;
  assign PE_109_reset = reset;
  assign PE_109_io_data_2_sig_stat2trans = PENetwork_56_io_to_pes_21_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_109_io_data_1_in_valid = PENetwork_26_io_to_pes_21_in_valid; // @[pe.scala 264:34]
  assign PE_109_io_data_1_in_bits = PENetwork_26_io_to_pes_21_in_bits; // @[pe.scala 264:34]
  assign PE_109_io_data_0_in_valid = PENetwork_21_io_to_pes_4_in_valid; // @[pe.scala 264:34]
  assign PE_109_io_data_0_in_bits = PENetwork_21_io_to_pes_4_in_bits; // @[pe.scala 264:34]
  assign PE_110_clock = clock;
  assign PE_110_reset = reset;
  assign PE_110_io_data_2_sig_stat2trans = PENetwork_57_io_to_pes_0_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_110_io_data_1_in_valid = PENetwork_27_io_to_pes_0_in_valid; // @[pe.scala 264:34]
  assign PE_110_io_data_1_in_bits = PENetwork_27_io_to_pes_0_in_bits; // @[pe.scala 264:34]
  assign PE_110_io_data_0_in_valid = PENetwork_io_to_pes_5_in_valid; // @[pe.scala 264:34]
  assign PE_110_io_data_0_in_bits = PENetwork_io_to_pes_5_in_bits; // @[pe.scala 264:34]
  assign PE_111_clock = clock;
  assign PE_111_reset = reset;
  assign PE_111_io_data_2_sig_stat2trans = PENetwork_57_io_to_pes_1_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_111_io_data_1_in_valid = PENetwork_27_io_to_pes_1_in_valid; // @[pe.scala 264:34]
  assign PE_111_io_data_1_in_bits = PENetwork_27_io_to_pes_1_in_bits; // @[pe.scala 264:34]
  assign PE_111_io_data_0_in_valid = PENetwork_1_io_to_pes_5_in_valid; // @[pe.scala 264:34]
  assign PE_111_io_data_0_in_bits = PENetwork_1_io_to_pes_5_in_bits; // @[pe.scala 264:34]
  assign PE_112_clock = clock;
  assign PE_112_reset = reset;
  assign PE_112_io_data_2_sig_stat2trans = PENetwork_57_io_to_pes_2_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_112_io_data_1_in_valid = PENetwork_27_io_to_pes_2_in_valid; // @[pe.scala 264:34]
  assign PE_112_io_data_1_in_bits = PENetwork_27_io_to_pes_2_in_bits; // @[pe.scala 264:34]
  assign PE_112_io_data_0_in_valid = PENetwork_2_io_to_pes_5_in_valid; // @[pe.scala 264:34]
  assign PE_112_io_data_0_in_bits = PENetwork_2_io_to_pes_5_in_bits; // @[pe.scala 264:34]
  assign PE_113_clock = clock;
  assign PE_113_reset = reset;
  assign PE_113_io_data_2_sig_stat2trans = PENetwork_57_io_to_pes_3_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_113_io_data_1_in_valid = PENetwork_27_io_to_pes_3_in_valid; // @[pe.scala 264:34]
  assign PE_113_io_data_1_in_bits = PENetwork_27_io_to_pes_3_in_bits; // @[pe.scala 264:34]
  assign PE_113_io_data_0_in_valid = PENetwork_3_io_to_pes_5_in_valid; // @[pe.scala 264:34]
  assign PE_113_io_data_0_in_bits = PENetwork_3_io_to_pes_5_in_bits; // @[pe.scala 264:34]
  assign PE_114_clock = clock;
  assign PE_114_reset = reset;
  assign PE_114_io_data_2_sig_stat2trans = PENetwork_57_io_to_pes_4_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_114_io_data_1_in_valid = PENetwork_27_io_to_pes_4_in_valid; // @[pe.scala 264:34]
  assign PE_114_io_data_1_in_bits = PENetwork_27_io_to_pes_4_in_bits; // @[pe.scala 264:34]
  assign PE_114_io_data_0_in_valid = PENetwork_4_io_to_pes_5_in_valid; // @[pe.scala 264:34]
  assign PE_114_io_data_0_in_bits = PENetwork_4_io_to_pes_5_in_bits; // @[pe.scala 264:34]
  assign PE_115_clock = clock;
  assign PE_115_reset = reset;
  assign PE_115_io_data_2_sig_stat2trans = PENetwork_57_io_to_pes_5_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_115_io_data_1_in_valid = PENetwork_27_io_to_pes_5_in_valid; // @[pe.scala 264:34]
  assign PE_115_io_data_1_in_bits = PENetwork_27_io_to_pes_5_in_bits; // @[pe.scala 264:34]
  assign PE_115_io_data_0_in_valid = PENetwork_5_io_to_pes_5_in_valid; // @[pe.scala 264:34]
  assign PE_115_io_data_0_in_bits = PENetwork_5_io_to_pes_5_in_bits; // @[pe.scala 264:34]
  assign PE_116_clock = clock;
  assign PE_116_reset = reset;
  assign PE_116_io_data_2_sig_stat2trans = PENetwork_57_io_to_pes_6_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_116_io_data_1_in_valid = PENetwork_27_io_to_pes_6_in_valid; // @[pe.scala 264:34]
  assign PE_116_io_data_1_in_bits = PENetwork_27_io_to_pes_6_in_bits; // @[pe.scala 264:34]
  assign PE_116_io_data_0_in_valid = PENetwork_6_io_to_pes_5_in_valid; // @[pe.scala 264:34]
  assign PE_116_io_data_0_in_bits = PENetwork_6_io_to_pes_5_in_bits; // @[pe.scala 264:34]
  assign PE_117_clock = clock;
  assign PE_117_reset = reset;
  assign PE_117_io_data_2_sig_stat2trans = PENetwork_57_io_to_pes_7_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_117_io_data_1_in_valid = PENetwork_27_io_to_pes_7_in_valid; // @[pe.scala 264:34]
  assign PE_117_io_data_1_in_bits = PENetwork_27_io_to_pes_7_in_bits; // @[pe.scala 264:34]
  assign PE_117_io_data_0_in_valid = PENetwork_7_io_to_pes_5_in_valid; // @[pe.scala 264:34]
  assign PE_117_io_data_0_in_bits = PENetwork_7_io_to_pes_5_in_bits; // @[pe.scala 264:34]
  assign PE_118_clock = clock;
  assign PE_118_reset = reset;
  assign PE_118_io_data_2_sig_stat2trans = PENetwork_57_io_to_pes_8_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_118_io_data_1_in_valid = PENetwork_27_io_to_pes_8_in_valid; // @[pe.scala 264:34]
  assign PE_118_io_data_1_in_bits = PENetwork_27_io_to_pes_8_in_bits; // @[pe.scala 264:34]
  assign PE_118_io_data_0_in_valid = PENetwork_8_io_to_pes_5_in_valid; // @[pe.scala 264:34]
  assign PE_118_io_data_0_in_bits = PENetwork_8_io_to_pes_5_in_bits; // @[pe.scala 264:34]
  assign PE_119_clock = clock;
  assign PE_119_reset = reset;
  assign PE_119_io_data_2_sig_stat2trans = PENetwork_57_io_to_pes_9_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_119_io_data_1_in_valid = PENetwork_27_io_to_pes_9_in_valid; // @[pe.scala 264:34]
  assign PE_119_io_data_1_in_bits = PENetwork_27_io_to_pes_9_in_bits; // @[pe.scala 264:34]
  assign PE_119_io_data_0_in_valid = PENetwork_9_io_to_pes_5_in_valid; // @[pe.scala 264:34]
  assign PE_119_io_data_0_in_bits = PENetwork_9_io_to_pes_5_in_bits; // @[pe.scala 264:34]
  assign PE_120_clock = clock;
  assign PE_120_reset = reset;
  assign PE_120_io_data_2_sig_stat2trans = PENetwork_57_io_to_pes_10_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_120_io_data_1_in_valid = PENetwork_27_io_to_pes_10_in_valid; // @[pe.scala 264:34]
  assign PE_120_io_data_1_in_bits = PENetwork_27_io_to_pes_10_in_bits; // @[pe.scala 264:34]
  assign PE_120_io_data_0_in_valid = PENetwork_10_io_to_pes_5_in_valid; // @[pe.scala 264:34]
  assign PE_120_io_data_0_in_bits = PENetwork_10_io_to_pes_5_in_bits; // @[pe.scala 264:34]
  assign PE_121_clock = clock;
  assign PE_121_reset = reset;
  assign PE_121_io_data_2_sig_stat2trans = PENetwork_57_io_to_pes_11_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_121_io_data_1_in_valid = PENetwork_27_io_to_pes_11_in_valid; // @[pe.scala 264:34]
  assign PE_121_io_data_1_in_bits = PENetwork_27_io_to_pes_11_in_bits; // @[pe.scala 264:34]
  assign PE_121_io_data_0_in_valid = PENetwork_11_io_to_pes_5_in_valid; // @[pe.scala 264:34]
  assign PE_121_io_data_0_in_bits = PENetwork_11_io_to_pes_5_in_bits; // @[pe.scala 264:34]
  assign PE_122_clock = clock;
  assign PE_122_reset = reset;
  assign PE_122_io_data_2_sig_stat2trans = PENetwork_57_io_to_pes_12_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_122_io_data_1_in_valid = PENetwork_27_io_to_pes_12_in_valid; // @[pe.scala 264:34]
  assign PE_122_io_data_1_in_bits = PENetwork_27_io_to_pes_12_in_bits; // @[pe.scala 264:34]
  assign PE_122_io_data_0_in_valid = PENetwork_12_io_to_pes_5_in_valid; // @[pe.scala 264:34]
  assign PE_122_io_data_0_in_bits = PENetwork_12_io_to_pes_5_in_bits; // @[pe.scala 264:34]
  assign PE_123_clock = clock;
  assign PE_123_reset = reset;
  assign PE_123_io_data_2_sig_stat2trans = PENetwork_57_io_to_pes_13_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_123_io_data_1_in_valid = PENetwork_27_io_to_pes_13_in_valid; // @[pe.scala 264:34]
  assign PE_123_io_data_1_in_bits = PENetwork_27_io_to_pes_13_in_bits; // @[pe.scala 264:34]
  assign PE_123_io_data_0_in_valid = PENetwork_13_io_to_pes_5_in_valid; // @[pe.scala 264:34]
  assign PE_123_io_data_0_in_bits = PENetwork_13_io_to_pes_5_in_bits; // @[pe.scala 264:34]
  assign PE_124_clock = clock;
  assign PE_124_reset = reset;
  assign PE_124_io_data_2_sig_stat2trans = PENetwork_57_io_to_pes_14_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_124_io_data_1_in_valid = PENetwork_27_io_to_pes_14_in_valid; // @[pe.scala 264:34]
  assign PE_124_io_data_1_in_bits = PENetwork_27_io_to_pes_14_in_bits; // @[pe.scala 264:34]
  assign PE_124_io_data_0_in_valid = PENetwork_14_io_to_pes_5_in_valid; // @[pe.scala 264:34]
  assign PE_124_io_data_0_in_bits = PENetwork_14_io_to_pes_5_in_bits; // @[pe.scala 264:34]
  assign PE_125_clock = clock;
  assign PE_125_reset = reset;
  assign PE_125_io_data_2_sig_stat2trans = PENetwork_57_io_to_pes_15_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_125_io_data_1_in_valid = PENetwork_27_io_to_pes_15_in_valid; // @[pe.scala 264:34]
  assign PE_125_io_data_1_in_bits = PENetwork_27_io_to_pes_15_in_bits; // @[pe.scala 264:34]
  assign PE_125_io_data_0_in_valid = PENetwork_15_io_to_pes_5_in_valid; // @[pe.scala 264:34]
  assign PE_125_io_data_0_in_bits = PENetwork_15_io_to_pes_5_in_bits; // @[pe.scala 264:34]
  assign PE_126_clock = clock;
  assign PE_126_reset = reset;
  assign PE_126_io_data_2_sig_stat2trans = PENetwork_57_io_to_pes_16_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_126_io_data_1_in_valid = PENetwork_27_io_to_pes_16_in_valid; // @[pe.scala 264:34]
  assign PE_126_io_data_1_in_bits = PENetwork_27_io_to_pes_16_in_bits; // @[pe.scala 264:34]
  assign PE_126_io_data_0_in_valid = PENetwork_16_io_to_pes_5_in_valid; // @[pe.scala 264:34]
  assign PE_126_io_data_0_in_bits = PENetwork_16_io_to_pes_5_in_bits; // @[pe.scala 264:34]
  assign PE_127_clock = clock;
  assign PE_127_reset = reset;
  assign PE_127_io_data_2_sig_stat2trans = PENetwork_57_io_to_pes_17_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_127_io_data_1_in_valid = PENetwork_27_io_to_pes_17_in_valid; // @[pe.scala 264:34]
  assign PE_127_io_data_1_in_bits = PENetwork_27_io_to_pes_17_in_bits; // @[pe.scala 264:34]
  assign PE_127_io_data_0_in_valid = PENetwork_17_io_to_pes_5_in_valid; // @[pe.scala 264:34]
  assign PE_127_io_data_0_in_bits = PENetwork_17_io_to_pes_5_in_bits; // @[pe.scala 264:34]
  assign PE_128_clock = clock;
  assign PE_128_reset = reset;
  assign PE_128_io_data_2_sig_stat2trans = PENetwork_57_io_to_pes_18_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_128_io_data_1_in_valid = PENetwork_27_io_to_pes_18_in_valid; // @[pe.scala 264:34]
  assign PE_128_io_data_1_in_bits = PENetwork_27_io_to_pes_18_in_bits; // @[pe.scala 264:34]
  assign PE_128_io_data_0_in_valid = PENetwork_18_io_to_pes_5_in_valid; // @[pe.scala 264:34]
  assign PE_128_io_data_0_in_bits = PENetwork_18_io_to_pes_5_in_bits; // @[pe.scala 264:34]
  assign PE_129_clock = clock;
  assign PE_129_reset = reset;
  assign PE_129_io_data_2_sig_stat2trans = PENetwork_57_io_to_pes_19_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_129_io_data_1_in_valid = PENetwork_27_io_to_pes_19_in_valid; // @[pe.scala 264:34]
  assign PE_129_io_data_1_in_bits = PENetwork_27_io_to_pes_19_in_bits; // @[pe.scala 264:34]
  assign PE_129_io_data_0_in_valid = PENetwork_19_io_to_pes_5_in_valid; // @[pe.scala 264:34]
  assign PE_129_io_data_0_in_bits = PENetwork_19_io_to_pes_5_in_bits; // @[pe.scala 264:34]
  assign PE_130_clock = clock;
  assign PE_130_reset = reset;
  assign PE_130_io_data_2_sig_stat2trans = PENetwork_57_io_to_pes_20_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_130_io_data_1_in_valid = PENetwork_27_io_to_pes_20_in_valid; // @[pe.scala 264:34]
  assign PE_130_io_data_1_in_bits = PENetwork_27_io_to_pes_20_in_bits; // @[pe.scala 264:34]
  assign PE_130_io_data_0_in_valid = PENetwork_20_io_to_pes_5_in_valid; // @[pe.scala 264:34]
  assign PE_130_io_data_0_in_bits = PENetwork_20_io_to_pes_5_in_bits; // @[pe.scala 264:34]
  assign PE_131_clock = clock;
  assign PE_131_reset = reset;
  assign PE_131_io_data_2_sig_stat2trans = PENetwork_57_io_to_pes_21_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_131_io_data_1_in_valid = PENetwork_27_io_to_pes_21_in_valid; // @[pe.scala 264:34]
  assign PE_131_io_data_1_in_bits = PENetwork_27_io_to_pes_21_in_bits; // @[pe.scala 264:34]
  assign PE_131_io_data_0_in_valid = PENetwork_21_io_to_pes_5_in_valid; // @[pe.scala 264:34]
  assign PE_131_io_data_0_in_bits = PENetwork_21_io_to_pes_5_in_bits; // @[pe.scala 264:34]
  assign PE_132_clock = clock;
  assign PE_132_reset = reset;
  assign PE_132_io_data_2_sig_stat2trans = PENetwork_58_io_to_pes_0_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_132_io_data_1_in_valid = PENetwork_28_io_to_pes_0_in_valid; // @[pe.scala 264:34]
  assign PE_132_io_data_1_in_bits = PENetwork_28_io_to_pes_0_in_bits; // @[pe.scala 264:34]
  assign PE_132_io_data_0_in_valid = PENetwork_io_to_pes_6_in_valid; // @[pe.scala 264:34]
  assign PE_132_io_data_0_in_bits = PENetwork_io_to_pes_6_in_bits; // @[pe.scala 264:34]
  assign PE_133_clock = clock;
  assign PE_133_reset = reset;
  assign PE_133_io_data_2_sig_stat2trans = PENetwork_58_io_to_pes_1_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_133_io_data_1_in_valid = PENetwork_28_io_to_pes_1_in_valid; // @[pe.scala 264:34]
  assign PE_133_io_data_1_in_bits = PENetwork_28_io_to_pes_1_in_bits; // @[pe.scala 264:34]
  assign PE_133_io_data_0_in_valid = PENetwork_1_io_to_pes_6_in_valid; // @[pe.scala 264:34]
  assign PE_133_io_data_0_in_bits = PENetwork_1_io_to_pes_6_in_bits; // @[pe.scala 264:34]
  assign PE_134_clock = clock;
  assign PE_134_reset = reset;
  assign PE_134_io_data_2_sig_stat2trans = PENetwork_58_io_to_pes_2_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_134_io_data_1_in_valid = PENetwork_28_io_to_pes_2_in_valid; // @[pe.scala 264:34]
  assign PE_134_io_data_1_in_bits = PENetwork_28_io_to_pes_2_in_bits; // @[pe.scala 264:34]
  assign PE_134_io_data_0_in_valid = PENetwork_2_io_to_pes_6_in_valid; // @[pe.scala 264:34]
  assign PE_134_io_data_0_in_bits = PENetwork_2_io_to_pes_6_in_bits; // @[pe.scala 264:34]
  assign PE_135_clock = clock;
  assign PE_135_reset = reset;
  assign PE_135_io_data_2_sig_stat2trans = PENetwork_58_io_to_pes_3_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_135_io_data_1_in_valid = PENetwork_28_io_to_pes_3_in_valid; // @[pe.scala 264:34]
  assign PE_135_io_data_1_in_bits = PENetwork_28_io_to_pes_3_in_bits; // @[pe.scala 264:34]
  assign PE_135_io_data_0_in_valid = PENetwork_3_io_to_pes_6_in_valid; // @[pe.scala 264:34]
  assign PE_135_io_data_0_in_bits = PENetwork_3_io_to_pes_6_in_bits; // @[pe.scala 264:34]
  assign PE_136_clock = clock;
  assign PE_136_reset = reset;
  assign PE_136_io_data_2_sig_stat2trans = PENetwork_58_io_to_pes_4_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_136_io_data_1_in_valid = PENetwork_28_io_to_pes_4_in_valid; // @[pe.scala 264:34]
  assign PE_136_io_data_1_in_bits = PENetwork_28_io_to_pes_4_in_bits; // @[pe.scala 264:34]
  assign PE_136_io_data_0_in_valid = PENetwork_4_io_to_pes_6_in_valid; // @[pe.scala 264:34]
  assign PE_136_io_data_0_in_bits = PENetwork_4_io_to_pes_6_in_bits; // @[pe.scala 264:34]
  assign PE_137_clock = clock;
  assign PE_137_reset = reset;
  assign PE_137_io_data_2_sig_stat2trans = PENetwork_58_io_to_pes_5_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_137_io_data_1_in_valid = PENetwork_28_io_to_pes_5_in_valid; // @[pe.scala 264:34]
  assign PE_137_io_data_1_in_bits = PENetwork_28_io_to_pes_5_in_bits; // @[pe.scala 264:34]
  assign PE_137_io_data_0_in_valid = PENetwork_5_io_to_pes_6_in_valid; // @[pe.scala 264:34]
  assign PE_137_io_data_0_in_bits = PENetwork_5_io_to_pes_6_in_bits; // @[pe.scala 264:34]
  assign PE_138_clock = clock;
  assign PE_138_reset = reset;
  assign PE_138_io_data_2_sig_stat2trans = PENetwork_58_io_to_pes_6_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_138_io_data_1_in_valid = PENetwork_28_io_to_pes_6_in_valid; // @[pe.scala 264:34]
  assign PE_138_io_data_1_in_bits = PENetwork_28_io_to_pes_6_in_bits; // @[pe.scala 264:34]
  assign PE_138_io_data_0_in_valid = PENetwork_6_io_to_pes_6_in_valid; // @[pe.scala 264:34]
  assign PE_138_io_data_0_in_bits = PENetwork_6_io_to_pes_6_in_bits; // @[pe.scala 264:34]
  assign PE_139_clock = clock;
  assign PE_139_reset = reset;
  assign PE_139_io_data_2_sig_stat2trans = PENetwork_58_io_to_pes_7_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_139_io_data_1_in_valid = PENetwork_28_io_to_pes_7_in_valid; // @[pe.scala 264:34]
  assign PE_139_io_data_1_in_bits = PENetwork_28_io_to_pes_7_in_bits; // @[pe.scala 264:34]
  assign PE_139_io_data_0_in_valid = PENetwork_7_io_to_pes_6_in_valid; // @[pe.scala 264:34]
  assign PE_139_io_data_0_in_bits = PENetwork_7_io_to_pes_6_in_bits; // @[pe.scala 264:34]
  assign PE_140_clock = clock;
  assign PE_140_reset = reset;
  assign PE_140_io_data_2_sig_stat2trans = PENetwork_58_io_to_pes_8_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_140_io_data_1_in_valid = PENetwork_28_io_to_pes_8_in_valid; // @[pe.scala 264:34]
  assign PE_140_io_data_1_in_bits = PENetwork_28_io_to_pes_8_in_bits; // @[pe.scala 264:34]
  assign PE_140_io_data_0_in_valid = PENetwork_8_io_to_pes_6_in_valid; // @[pe.scala 264:34]
  assign PE_140_io_data_0_in_bits = PENetwork_8_io_to_pes_6_in_bits; // @[pe.scala 264:34]
  assign PE_141_clock = clock;
  assign PE_141_reset = reset;
  assign PE_141_io_data_2_sig_stat2trans = PENetwork_58_io_to_pes_9_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_141_io_data_1_in_valid = PENetwork_28_io_to_pes_9_in_valid; // @[pe.scala 264:34]
  assign PE_141_io_data_1_in_bits = PENetwork_28_io_to_pes_9_in_bits; // @[pe.scala 264:34]
  assign PE_141_io_data_0_in_valid = PENetwork_9_io_to_pes_6_in_valid; // @[pe.scala 264:34]
  assign PE_141_io_data_0_in_bits = PENetwork_9_io_to_pes_6_in_bits; // @[pe.scala 264:34]
  assign PE_142_clock = clock;
  assign PE_142_reset = reset;
  assign PE_142_io_data_2_sig_stat2trans = PENetwork_58_io_to_pes_10_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_142_io_data_1_in_valid = PENetwork_28_io_to_pes_10_in_valid; // @[pe.scala 264:34]
  assign PE_142_io_data_1_in_bits = PENetwork_28_io_to_pes_10_in_bits; // @[pe.scala 264:34]
  assign PE_142_io_data_0_in_valid = PENetwork_10_io_to_pes_6_in_valid; // @[pe.scala 264:34]
  assign PE_142_io_data_0_in_bits = PENetwork_10_io_to_pes_6_in_bits; // @[pe.scala 264:34]
  assign PE_143_clock = clock;
  assign PE_143_reset = reset;
  assign PE_143_io_data_2_sig_stat2trans = PENetwork_58_io_to_pes_11_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_143_io_data_1_in_valid = PENetwork_28_io_to_pes_11_in_valid; // @[pe.scala 264:34]
  assign PE_143_io_data_1_in_bits = PENetwork_28_io_to_pes_11_in_bits; // @[pe.scala 264:34]
  assign PE_143_io_data_0_in_valid = PENetwork_11_io_to_pes_6_in_valid; // @[pe.scala 264:34]
  assign PE_143_io_data_0_in_bits = PENetwork_11_io_to_pes_6_in_bits; // @[pe.scala 264:34]
  assign PE_144_clock = clock;
  assign PE_144_reset = reset;
  assign PE_144_io_data_2_sig_stat2trans = PENetwork_58_io_to_pes_12_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_144_io_data_1_in_valid = PENetwork_28_io_to_pes_12_in_valid; // @[pe.scala 264:34]
  assign PE_144_io_data_1_in_bits = PENetwork_28_io_to_pes_12_in_bits; // @[pe.scala 264:34]
  assign PE_144_io_data_0_in_valid = PENetwork_12_io_to_pes_6_in_valid; // @[pe.scala 264:34]
  assign PE_144_io_data_0_in_bits = PENetwork_12_io_to_pes_6_in_bits; // @[pe.scala 264:34]
  assign PE_145_clock = clock;
  assign PE_145_reset = reset;
  assign PE_145_io_data_2_sig_stat2trans = PENetwork_58_io_to_pes_13_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_145_io_data_1_in_valid = PENetwork_28_io_to_pes_13_in_valid; // @[pe.scala 264:34]
  assign PE_145_io_data_1_in_bits = PENetwork_28_io_to_pes_13_in_bits; // @[pe.scala 264:34]
  assign PE_145_io_data_0_in_valid = PENetwork_13_io_to_pes_6_in_valid; // @[pe.scala 264:34]
  assign PE_145_io_data_0_in_bits = PENetwork_13_io_to_pes_6_in_bits; // @[pe.scala 264:34]
  assign PE_146_clock = clock;
  assign PE_146_reset = reset;
  assign PE_146_io_data_2_sig_stat2trans = PENetwork_58_io_to_pes_14_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_146_io_data_1_in_valid = PENetwork_28_io_to_pes_14_in_valid; // @[pe.scala 264:34]
  assign PE_146_io_data_1_in_bits = PENetwork_28_io_to_pes_14_in_bits; // @[pe.scala 264:34]
  assign PE_146_io_data_0_in_valid = PENetwork_14_io_to_pes_6_in_valid; // @[pe.scala 264:34]
  assign PE_146_io_data_0_in_bits = PENetwork_14_io_to_pes_6_in_bits; // @[pe.scala 264:34]
  assign PE_147_clock = clock;
  assign PE_147_reset = reset;
  assign PE_147_io_data_2_sig_stat2trans = PENetwork_58_io_to_pes_15_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_147_io_data_1_in_valid = PENetwork_28_io_to_pes_15_in_valid; // @[pe.scala 264:34]
  assign PE_147_io_data_1_in_bits = PENetwork_28_io_to_pes_15_in_bits; // @[pe.scala 264:34]
  assign PE_147_io_data_0_in_valid = PENetwork_15_io_to_pes_6_in_valid; // @[pe.scala 264:34]
  assign PE_147_io_data_0_in_bits = PENetwork_15_io_to_pes_6_in_bits; // @[pe.scala 264:34]
  assign PE_148_clock = clock;
  assign PE_148_reset = reset;
  assign PE_148_io_data_2_sig_stat2trans = PENetwork_58_io_to_pes_16_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_148_io_data_1_in_valid = PENetwork_28_io_to_pes_16_in_valid; // @[pe.scala 264:34]
  assign PE_148_io_data_1_in_bits = PENetwork_28_io_to_pes_16_in_bits; // @[pe.scala 264:34]
  assign PE_148_io_data_0_in_valid = PENetwork_16_io_to_pes_6_in_valid; // @[pe.scala 264:34]
  assign PE_148_io_data_0_in_bits = PENetwork_16_io_to_pes_6_in_bits; // @[pe.scala 264:34]
  assign PE_149_clock = clock;
  assign PE_149_reset = reset;
  assign PE_149_io_data_2_sig_stat2trans = PENetwork_58_io_to_pes_17_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_149_io_data_1_in_valid = PENetwork_28_io_to_pes_17_in_valid; // @[pe.scala 264:34]
  assign PE_149_io_data_1_in_bits = PENetwork_28_io_to_pes_17_in_bits; // @[pe.scala 264:34]
  assign PE_149_io_data_0_in_valid = PENetwork_17_io_to_pes_6_in_valid; // @[pe.scala 264:34]
  assign PE_149_io_data_0_in_bits = PENetwork_17_io_to_pes_6_in_bits; // @[pe.scala 264:34]
  assign PE_150_clock = clock;
  assign PE_150_reset = reset;
  assign PE_150_io_data_2_sig_stat2trans = PENetwork_58_io_to_pes_18_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_150_io_data_1_in_valid = PENetwork_28_io_to_pes_18_in_valid; // @[pe.scala 264:34]
  assign PE_150_io_data_1_in_bits = PENetwork_28_io_to_pes_18_in_bits; // @[pe.scala 264:34]
  assign PE_150_io_data_0_in_valid = PENetwork_18_io_to_pes_6_in_valid; // @[pe.scala 264:34]
  assign PE_150_io_data_0_in_bits = PENetwork_18_io_to_pes_6_in_bits; // @[pe.scala 264:34]
  assign PE_151_clock = clock;
  assign PE_151_reset = reset;
  assign PE_151_io_data_2_sig_stat2trans = PENetwork_58_io_to_pes_19_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_151_io_data_1_in_valid = PENetwork_28_io_to_pes_19_in_valid; // @[pe.scala 264:34]
  assign PE_151_io_data_1_in_bits = PENetwork_28_io_to_pes_19_in_bits; // @[pe.scala 264:34]
  assign PE_151_io_data_0_in_valid = PENetwork_19_io_to_pes_6_in_valid; // @[pe.scala 264:34]
  assign PE_151_io_data_0_in_bits = PENetwork_19_io_to_pes_6_in_bits; // @[pe.scala 264:34]
  assign PE_152_clock = clock;
  assign PE_152_reset = reset;
  assign PE_152_io_data_2_sig_stat2trans = PENetwork_58_io_to_pes_20_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_152_io_data_1_in_valid = PENetwork_28_io_to_pes_20_in_valid; // @[pe.scala 264:34]
  assign PE_152_io_data_1_in_bits = PENetwork_28_io_to_pes_20_in_bits; // @[pe.scala 264:34]
  assign PE_152_io_data_0_in_valid = PENetwork_20_io_to_pes_6_in_valid; // @[pe.scala 264:34]
  assign PE_152_io_data_0_in_bits = PENetwork_20_io_to_pes_6_in_bits; // @[pe.scala 264:34]
  assign PE_153_clock = clock;
  assign PE_153_reset = reset;
  assign PE_153_io_data_2_sig_stat2trans = PENetwork_58_io_to_pes_21_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_153_io_data_1_in_valid = PENetwork_28_io_to_pes_21_in_valid; // @[pe.scala 264:34]
  assign PE_153_io_data_1_in_bits = PENetwork_28_io_to_pes_21_in_bits; // @[pe.scala 264:34]
  assign PE_153_io_data_0_in_valid = PENetwork_21_io_to_pes_6_in_valid; // @[pe.scala 264:34]
  assign PE_153_io_data_0_in_bits = PENetwork_21_io_to_pes_6_in_bits; // @[pe.scala 264:34]
  assign PE_154_clock = clock;
  assign PE_154_reset = reset;
  assign PE_154_io_data_2_sig_stat2trans = PENetwork_59_io_to_pes_0_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_154_io_data_1_in_valid = PENetwork_29_io_to_pes_0_in_valid; // @[pe.scala 264:34]
  assign PE_154_io_data_1_in_bits = PENetwork_29_io_to_pes_0_in_bits; // @[pe.scala 264:34]
  assign PE_154_io_data_0_in_valid = PENetwork_io_to_pes_7_in_valid; // @[pe.scala 264:34]
  assign PE_154_io_data_0_in_bits = PENetwork_io_to_pes_7_in_bits; // @[pe.scala 264:34]
  assign PE_155_clock = clock;
  assign PE_155_reset = reset;
  assign PE_155_io_data_2_sig_stat2trans = PENetwork_59_io_to_pes_1_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_155_io_data_1_in_valid = PENetwork_29_io_to_pes_1_in_valid; // @[pe.scala 264:34]
  assign PE_155_io_data_1_in_bits = PENetwork_29_io_to_pes_1_in_bits; // @[pe.scala 264:34]
  assign PE_155_io_data_0_in_valid = PENetwork_1_io_to_pes_7_in_valid; // @[pe.scala 264:34]
  assign PE_155_io_data_0_in_bits = PENetwork_1_io_to_pes_7_in_bits; // @[pe.scala 264:34]
  assign PE_156_clock = clock;
  assign PE_156_reset = reset;
  assign PE_156_io_data_2_sig_stat2trans = PENetwork_59_io_to_pes_2_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_156_io_data_1_in_valid = PENetwork_29_io_to_pes_2_in_valid; // @[pe.scala 264:34]
  assign PE_156_io_data_1_in_bits = PENetwork_29_io_to_pes_2_in_bits; // @[pe.scala 264:34]
  assign PE_156_io_data_0_in_valid = PENetwork_2_io_to_pes_7_in_valid; // @[pe.scala 264:34]
  assign PE_156_io_data_0_in_bits = PENetwork_2_io_to_pes_7_in_bits; // @[pe.scala 264:34]
  assign PE_157_clock = clock;
  assign PE_157_reset = reset;
  assign PE_157_io_data_2_sig_stat2trans = PENetwork_59_io_to_pes_3_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_157_io_data_1_in_valid = PENetwork_29_io_to_pes_3_in_valid; // @[pe.scala 264:34]
  assign PE_157_io_data_1_in_bits = PENetwork_29_io_to_pes_3_in_bits; // @[pe.scala 264:34]
  assign PE_157_io_data_0_in_valid = PENetwork_3_io_to_pes_7_in_valid; // @[pe.scala 264:34]
  assign PE_157_io_data_0_in_bits = PENetwork_3_io_to_pes_7_in_bits; // @[pe.scala 264:34]
  assign PE_158_clock = clock;
  assign PE_158_reset = reset;
  assign PE_158_io_data_2_sig_stat2trans = PENetwork_59_io_to_pes_4_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_158_io_data_1_in_valid = PENetwork_29_io_to_pes_4_in_valid; // @[pe.scala 264:34]
  assign PE_158_io_data_1_in_bits = PENetwork_29_io_to_pes_4_in_bits; // @[pe.scala 264:34]
  assign PE_158_io_data_0_in_valid = PENetwork_4_io_to_pes_7_in_valid; // @[pe.scala 264:34]
  assign PE_158_io_data_0_in_bits = PENetwork_4_io_to_pes_7_in_bits; // @[pe.scala 264:34]
  assign PE_159_clock = clock;
  assign PE_159_reset = reset;
  assign PE_159_io_data_2_sig_stat2trans = PENetwork_59_io_to_pes_5_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_159_io_data_1_in_valid = PENetwork_29_io_to_pes_5_in_valid; // @[pe.scala 264:34]
  assign PE_159_io_data_1_in_bits = PENetwork_29_io_to_pes_5_in_bits; // @[pe.scala 264:34]
  assign PE_159_io_data_0_in_valid = PENetwork_5_io_to_pes_7_in_valid; // @[pe.scala 264:34]
  assign PE_159_io_data_0_in_bits = PENetwork_5_io_to_pes_7_in_bits; // @[pe.scala 264:34]
  assign PE_160_clock = clock;
  assign PE_160_reset = reset;
  assign PE_160_io_data_2_sig_stat2trans = PENetwork_59_io_to_pes_6_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_160_io_data_1_in_valid = PENetwork_29_io_to_pes_6_in_valid; // @[pe.scala 264:34]
  assign PE_160_io_data_1_in_bits = PENetwork_29_io_to_pes_6_in_bits; // @[pe.scala 264:34]
  assign PE_160_io_data_0_in_valid = PENetwork_6_io_to_pes_7_in_valid; // @[pe.scala 264:34]
  assign PE_160_io_data_0_in_bits = PENetwork_6_io_to_pes_7_in_bits; // @[pe.scala 264:34]
  assign PE_161_clock = clock;
  assign PE_161_reset = reset;
  assign PE_161_io_data_2_sig_stat2trans = PENetwork_59_io_to_pes_7_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_161_io_data_1_in_valid = PENetwork_29_io_to_pes_7_in_valid; // @[pe.scala 264:34]
  assign PE_161_io_data_1_in_bits = PENetwork_29_io_to_pes_7_in_bits; // @[pe.scala 264:34]
  assign PE_161_io_data_0_in_valid = PENetwork_7_io_to_pes_7_in_valid; // @[pe.scala 264:34]
  assign PE_161_io_data_0_in_bits = PENetwork_7_io_to_pes_7_in_bits; // @[pe.scala 264:34]
  assign PE_162_clock = clock;
  assign PE_162_reset = reset;
  assign PE_162_io_data_2_sig_stat2trans = PENetwork_59_io_to_pes_8_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_162_io_data_1_in_valid = PENetwork_29_io_to_pes_8_in_valid; // @[pe.scala 264:34]
  assign PE_162_io_data_1_in_bits = PENetwork_29_io_to_pes_8_in_bits; // @[pe.scala 264:34]
  assign PE_162_io_data_0_in_valid = PENetwork_8_io_to_pes_7_in_valid; // @[pe.scala 264:34]
  assign PE_162_io_data_0_in_bits = PENetwork_8_io_to_pes_7_in_bits; // @[pe.scala 264:34]
  assign PE_163_clock = clock;
  assign PE_163_reset = reset;
  assign PE_163_io_data_2_sig_stat2trans = PENetwork_59_io_to_pes_9_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_163_io_data_1_in_valid = PENetwork_29_io_to_pes_9_in_valid; // @[pe.scala 264:34]
  assign PE_163_io_data_1_in_bits = PENetwork_29_io_to_pes_9_in_bits; // @[pe.scala 264:34]
  assign PE_163_io_data_0_in_valid = PENetwork_9_io_to_pes_7_in_valid; // @[pe.scala 264:34]
  assign PE_163_io_data_0_in_bits = PENetwork_9_io_to_pes_7_in_bits; // @[pe.scala 264:34]
  assign PE_164_clock = clock;
  assign PE_164_reset = reset;
  assign PE_164_io_data_2_sig_stat2trans = PENetwork_59_io_to_pes_10_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_164_io_data_1_in_valid = PENetwork_29_io_to_pes_10_in_valid; // @[pe.scala 264:34]
  assign PE_164_io_data_1_in_bits = PENetwork_29_io_to_pes_10_in_bits; // @[pe.scala 264:34]
  assign PE_164_io_data_0_in_valid = PENetwork_10_io_to_pes_7_in_valid; // @[pe.scala 264:34]
  assign PE_164_io_data_0_in_bits = PENetwork_10_io_to_pes_7_in_bits; // @[pe.scala 264:34]
  assign PE_165_clock = clock;
  assign PE_165_reset = reset;
  assign PE_165_io_data_2_sig_stat2trans = PENetwork_59_io_to_pes_11_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_165_io_data_1_in_valid = PENetwork_29_io_to_pes_11_in_valid; // @[pe.scala 264:34]
  assign PE_165_io_data_1_in_bits = PENetwork_29_io_to_pes_11_in_bits; // @[pe.scala 264:34]
  assign PE_165_io_data_0_in_valid = PENetwork_11_io_to_pes_7_in_valid; // @[pe.scala 264:34]
  assign PE_165_io_data_0_in_bits = PENetwork_11_io_to_pes_7_in_bits; // @[pe.scala 264:34]
  assign PE_166_clock = clock;
  assign PE_166_reset = reset;
  assign PE_166_io_data_2_sig_stat2trans = PENetwork_59_io_to_pes_12_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_166_io_data_1_in_valid = PENetwork_29_io_to_pes_12_in_valid; // @[pe.scala 264:34]
  assign PE_166_io_data_1_in_bits = PENetwork_29_io_to_pes_12_in_bits; // @[pe.scala 264:34]
  assign PE_166_io_data_0_in_valid = PENetwork_12_io_to_pes_7_in_valid; // @[pe.scala 264:34]
  assign PE_166_io_data_0_in_bits = PENetwork_12_io_to_pes_7_in_bits; // @[pe.scala 264:34]
  assign PE_167_clock = clock;
  assign PE_167_reset = reset;
  assign PE_167_io_data_2_sig_stat2trans = PENetwork_59_io_to_pes_13_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_167_io_data_1_in_valid = PENetwork_29_io_to_pes_13_in_valid; // @[pe.scala 264:34]
  assign PE_167_io_data_1_in_bits = PENetwork_29_io_to_pes_13_in_bits; // @[pe.scala 264:34]
  assign PE_167_io_data_0_in_valid = PENetwork_13_io_to_pes_7_in_valid; // @[pe.scala 264:34]
  assign PE_167_io_data_0_in_bits = PENetwork_13_io_to_pes_7_in_bits; // @[pe.scala 264:34]
  assign PE_168_clock = clock;
  assign PE_168_reset = reset;
  assign PE_168_io_data_2_sig_stat2trans = PENetwork_59_io_to_pes_14_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_168_io_data_1_in_valid = PENetwork_29_io_to_pes_14_in_valid; // @[pe.scala 264:34]
  assign PE_168_io_data_1_in_bits = PENetwork_29_io_to_pes_14_in_bits; // @[pe.scala 264:34]
  assign PE_168_io_data_0_in_valid = PENetwork_14_io_to_pes_7_in_valid; // @[pe.scala 264:34]
  assign PE_168_io_data_0_in_bits = PENetwork_14_io_to_pes_7_in_bits; // @[pe.scala 264:34]
  assign PE_169_clock = clock;
  assign PE_169_reset = reset;
  assign PE_169_io_data_2_sig_stat2trans = PENetwork_59_io_to_pes_15_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_169_io_data_1_in_valid = PENetwork_29_io_to_pes_15_in_valid; // @[pe.scala 264:34]
  assign PE_169_io_data_1_in_bits = PENetwork_29_io_to_pes_15_in_bits; // @[pe.scala 264:34]
  assign PE_169_io_data_0_in_valid = PENetwork_15_io_to_pes_7_in_valid; // @[pe.scala 264:34]
  assign PE_169_io_data_0_in_bits = PENetwork_15_io_to_pes_7_in_bits; // @[pe.scala 264:34]
  assign PE_170_clock = clock;
  assign PE_170_reset = reset;
  assign PE_170_io_data_2_sig_stat2trans = PENetwork_59_io_to_pes_16_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_170_io_data_1_in_valid = PENetwork_29_io_to_pes_16_in_valid; // @[pe.scala 264:34]
  assign PE_170_io_data_1_in_bits = PENetwork_29_io_to_pes_16_in_bits; // @[pe.scala 264:34]
  assign PE_170_io_data_0_in_valid = PENetwork_16_io_to_pes_7_in_valid; // @[pe.scala 264:34]
  assign PE_170_io_data_0_in_bits = PENetwork_16_io_to_pes_7_in_bits; // @[pe.scala 264:34]
  assign PE_171_clock = clock;
  assign PE_171_reset = reset;
  assign PE_171_io_data_2_sig_stat2trans = PENetwork_59_io_to_pes_17_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_171_io_data_1_in_valid = PENetwork_29_io_to_pes_17_in_valid; // @[pe.scala 264:34]
  assign PE_171_io_data_1_in_bits = PENetwork_29_io_to_pes_17_in_bits; // @[pe.scala 264:34]
  assign PE_171_io_data_0_in_valid = PENetwork_17_io_to_pes_7_in_valid; // @[pe.scala 264:34]
  assign PE_171_io_data_0_in_bits = PENetwork_17_io_to_pes_7_in_bits; // @[pe.scala 264:34]
  assign PE_172_clock = clock;
  assign PE_172_reset = reset;
  assign PE_172_io_data_2_sig_stat2trans = PENetwork_59_io_to_pes_18_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_172_io_data_1_in_valid = PENetwork_29_io_to_pes_18_in_valid; // @[pe.scala 264:34]
  assign PE_172_io_data_1_in_bits = PENetwork_29_io_to_pes_18_in_bits; // @[pe.scala 264:34]
  assign PE_172_io_data_0_in_valid = PENetwork_18_io_to_pes_7_in_valid; // @[pe.scala 264:34]
  assign PE_172_io_data_0_in_bits = PENetwork_18_io_to_pes_7_in_bits; // @[pe.scala 264:34]
  assign PE_173_clock = clock;
  assign PE_173_reset = reset;
  assign PE_173_io_data_2_sig_stat2trans = PENetwork_59_io_to_pes_19_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_173_io_data_1_in_valid = PENetwork_29_io_to_pes_19_in_valid; // @[pe.scala 264:34]
  assign PE_173_io_data_1_in_bits = PENetwork_29_io_to_pes_19_in_bits; // @[pe.scala 264:34]
  assign PE_173_io_data_0_in_valid = PENetwork_19_io_to_pes_7_in_valid; // @[pe.scala 264:34]
  assign PE_173_io_data_0_in_bits = PENetwork_19_io_to_pes_7_in_bits; // @[pe.scala 264:34]
  assign PE_174_clock = clock;
  assign PE_174_reset = reset;
  assign PE_174_io_data_2_sig_stat2trans = PENetwork_59_io_to_pes_20_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_174_io_data_1_in_valid = PENetwork_29_io_to_pes_20_in_valid; // @[pe.scala 264:34]
  assign PE_174_io_data_1_in_bits = PENetwork_29_io_to_pes_20_in_bits; // @[pe.scala 264:34]
  assign PE_174_io_data_0_in_valid = PENetwork_20_io_to_pes_7_in_valid; // @[pe.scala 264:34]
  assign PE_174_io_data_0_in_bits = PENetwork_20_io_to_pes_7_in_bits; // @[pe.scala 264:34]
  assign PE_175_clock = clock;
  assign PE_175_reset = reset;
  assign PE_175_io_data_2_sig_stat2trans = PENetwork_59_io_to_pes_21_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_175_io_data_1_in_valid = PENetwork_29_io_to_pes_21_in_valid; // @[pe.scala 264:34]
  assign PE_175_io_data_1_in_bits = PENetwork_29_io_to_pes_21_in_bits; // @[pe.scala 264:34]
  assign PE_175_io_data_0_in_valid = PENetwork_21_io_to_pes_7_in_valid; // @[pe.scala 264:34]
  assign PE_175_io_data_0_in_bits = PENetwork_21_io_to_pes_7_in_bits; // @[pe.scala 264:34]
  assign PE_176_clock = clock;
  assign PE_176_reset = reset;
  assign PE_176_io_data_2_sig_stat2trans = PENetwork_60_io_to_pes_0_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_176_io_data_1_in_valid = PENetwork_30_io_to_pes_0_in_valid; // @[pe.scala 264:34]
  assign PE_176_io_data_1_in_bits = PENetwork_30_io_to_pes_0_in_bits; // @[pe.scala 264:34]
  assign PE_176_io_data_0_in_valid = PENetwork_io_to_pes_8_in_valid; // @[pe.scala 264:34]
  assign PE_176_io_data_0_in_bits = PENetwork_io_to_pes_8_in_bits; // @[pe.scala 264:34]
  assign PE_177_clock = clock;
  assign PE_177_reset = reset;
  assign PE_177_io_data_2_sig_stat2trans = PENetwork_60_io_to_pes_1_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_177_io_data_1_in_valid = PENetwork_30_io_to_pes_1_in_valid; // @[pe.scala 264:34]
  assign PE_177_io_data_1_in_bits = PENetwork_30_io_to_pes_1_in_bits; // @[pe.scala 264:34]
  assign PE_177_io_data_0_in_valid = PENetwork_1_io_to_pes_8_in_valid; // @[pe.scala 264:34]
  assign PE_177_io_data_0_in_bits = PENetwork_1_io_to_pes_8_in_bits; // @[pe.scala 264:34]
  assign PE_178_clock = clock;
  assign PE_178_reset = reset;
  assign PE_178_io_data_2_sig_stat2trans = PENetwork_60_io_to_pes_2_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_178_io_data_1_in_valid = PENetwork_30_io_to_pes_2_in_valid; // @[pe.scala 264:34]
  assign PE_178_io_data_1_in_bits = PENetwork_30_io_to_pes_2_in_bits; // @[pe.scala 264:34]
  assign PE_178_io_data_0_in_valid = PENetwork_2_io_to_pes_8_in_valid; // @[pe.scala 264:34]
  assign PE_178_io_data_0_in_bits = PENetwork_2_io_to_pes_8_in_bits; // @[pe.scala 264:34]
  assign PE_179_clock = clock;
  assign PE_179_reset = reset;
  assign PE_179_io_data_2_sig_stat2trans = PENetwork_60_io_to_pes_3_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_179_io_data_1_in_valid = PENetwork_30_io_to_pes_3_in_valid; // @[pe.scala 264:34]
  assign PE_179_io_data_1_in_bits = PENetwork_30_io_to_pes_3_in_bits; // @[pe.scala 264:34]
  assign PE_179_io_data_0_in_valid = PENetwork_3_io_to_pes_8_in_valid; // @[pe.scala 264:34]
  assign PE_179_io_data_0_in_bits = PENetwork_3_io_to_pes_8_in_bits; // @[pe.scala 264:34]
  assign PE_180_clock = clock;
  assign PE_180_reset = reset;
  assign PE_180_io_data_2_sig_stat2trans = PENetwork_60_io_to_pes_4_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_180_io_data_1_in_valid = PENetwork_30_io_to_pes_4_in_valid; // @[pe.scala 264:34]
  assign PE_180_io_data_1_in_bits = PENetwork_30_io_to_pes_4_in_bits; // @[pe.scala 264:34]
  assign PE_180_io_data_0_in_valid = PENetwork_4_io_to_pes_8_in_valid; // @[pe.scala 264:34]
  assign PE_180_io_data_0_in_bits = PENetwork_4_io_to_pes_8_in_bits; // @[pe.scala 264:34]
  assign PE_181_clock = clock;
  assign PE_181_reset = reset;
  assign PE_181_io_data_2_sig_stat2trans = PENetwork_60_io_to_pes_5_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_181_io_data_1_in_valid = PENetwork_30_io_to_pes_5_in_valid; // @[pe.scala 264:34]
  assign PE_181_io_data_1_in_bits = PENetwork_30_io_to_pes_5_in_bits; // @[pe.scala 264:34]
  assign PE_181_io_data_0_in_valid = PENetwork_5_io_to_pes_8_in_valid; // @[pe.scala 264:34]
  assign PE_181_io_data_0_in_bits = PENetwork_5_io_to_pes_8_in_bits; // @[pe.scala 264:34]
  assign PE_182_clock = clock;
  assign PE_182_reset = reset;
  assign PE_182_io_data_2_sig_stat2trans = PENetwork_60_io_to_pes_6_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_182_io_data_1_in_valid = PENetwork_30_io_to_pes_6_in_valid; // @[pe.scala 264:34]
  assign PE_182_io_data_1_in_bits = PENetwork_30_io_to_pes_6_in_bits; // @[pe.scala 264:34]
  assign PE_182_io_data_0_in_valid = PENetwork_6_io_to_pes_8_in_valid; // @[pe.scala 264:34]
  assign PE_182_io_data_0_in_bits = PENetwork_6_io_to_pes_8_in_bits; // @[pe.scala 264:34]
  assign PE_183_clock = clock;
  assign PE_183_reset = reset;
  assign PE_183_io_data_2_sig_stat2trans = PENetwork_60_io_to_pes_7_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_183_io_data_1_in_valid = PENetwork_30_io_to_pes_7_in_valid; // @[pe.scala 264:34]
  assign PE_183_io_data_1_in_bits = PENetwork_30_io_to_pes_7_in_bits; // @[pe.scala 264:34]
  assign PE_183_io_data_0_in_valid = PENetwork_7_io_to_pes_8_in_valid; // @[pe.scala 264:34]
  assign PE_183_io_data_0_in_bits = PENetwork_7_io_to_pes_8_in_bits; // @[pe.scala 264:34]
  assign PE_184_clock = clock;
  assign PE_184_reset = reset;
  assign PE_184_io_data_2_sig_stat2trans = PENetwork_60_io_to_pes_8_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_184_io_data_1_in_valid = PENetwork_30_io_to_pes_8_in_valid; // @[pe.scala 264:34]
  assign PE_184_io_data_1_in_bits = PENetwork_30_io_to_pes_8_in_bits; // @[pe.scala 264:34]
  assign PE_184_io_data_0_in_valid = PENetwork_8_io_to_pes_8_in_valid; // @[pe.scala 264:34]
  assign PE_184_io_data_0_in_bits = PENetwork_8_io_to_pes_8_in_bits; // @[pe.scala 264:34]
  assign PE_185_clock = clock;
  assign PE_185_reset = reset;
  assign PE_185_io_data_2_sig_stat2trans = PENetwork_60_io_to_pes_9_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_185_io_data_1_in_valid = PENetwork_30_io_to_pes_9_in_valid; // @[pe.scala 264:34]
  assign PE_185_io_data_1_in_bits = PENetwork_30_io_to_pes_9_in_bits; // @[pe.scala 264:34]
  assign PE_185_io_data_0_in_valid = PENetwork_9_io_to_pes_8_in_valid; // @[pe.scala 264:34]
  assign PE_185_io_data_0_in_bits = PENetwork_9_io_to_pes_8_in_bits; // @[pe.scala 264:34]
  assign PE_186_clock = clock;
  assign PE_186_reset = reset;
  assign PE_186_io_data_2_sig_stat2trans = PENetwork_60_io_to_pes_10_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_186_io_data_1_in_valid = PENetwork_30_io_to_pes_10_in_valid; // @[pe.scala 264:34]
  assign PE_186_io_data_1_in_bits = PENetwork_30_io_to_pes_10_in_bits; // @[pe.scala 264:34]
  assign PE_186_io_data_0_in_valid = PENetwork_10_io_to_pes_8_in_valid; // @[pe.scala 264:34]
  assign PE_186_io_data_0_in_bits = PENetwork_10_io_to_pes_8_in_bits; // @[pe.scala 264:34]
  assign PE_187_clock = clock;
  assign PE_187_reset = reset;
  assign PE_187_io_data_2_sig_stat2trans = PENetwork_60_io_to_pes_11_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_187_io_data_1_in_valid = PENetwork_30_io_to_pes_11_in_valid; // @[pe.scala 264:34]
  assign PE_187_io_data_1_in_bits = PENetwork_30_io_to_pes_11_in_bits; // @[pe.scala 264:34]
  assign PE_187_io_data_0_in_valid = PENetwork_11_io_to_pes_8_in_valid; // @[pe.scala 264:34]
  assign PE_187_io_data_0_in_bits = PENetwork_11_io_to_pes_8_in_bits; // @[pe.scala 264:34]
  assign PE_188_clock = clock;
  assign PE_188_reset = reset;
  assign PE_188_io_data_2_sig_stat2trans = PENetwork_60_io_to_pes_12_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_188_io_data_1_in_valid = PENetwork_30_io_to_pes_12_in_valid; // @[pe.scala 264:34]
  assign PE_188_io_data_1_in_bits = PENetwork_30_io_to_pes_12_in_bits; // @[pe.scala 264:34]
  assign PE_188_io_data_0_in_valid = PENetwork_12_io_to_pes_8_in_valid; // @[pe.scala 264:34]
  assign PE_188_io_data_0_in_bits = PENetwork_12_io_to_pes_8_in_bits; // @[pe.scala 264:34]
  assign PE_189_clock = clock;
  assign PE_189_reset = reset;
  assign PE_189_io_data_2_sig_stat2trans = PENetwork_60_io_to_pes_13_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_189_io_data_1_in_valid = PENetwork_30_io_to_pes_13_in_valid; // @[pe.scala 264:34]
  assign PE_189_io_data_1_in_bits = PENetwork_30_io_to_pes_13_in_bits; // @[pe.scala 264:34]
  assign PE_189_io_data_0_in_valid = PENetwork_13_io_to_pes_8_in_valid; // @[pe.scala 264:34]
  assign PE_189_io_data_0_in_bits = PENetwork_13_io_to_pes_8_in_bits; // @[pe.scala 264:34]
  assign PE_190_clock = clock;
  assign PE_190_reset = reset;
  assign PE_190_io_data_2_sig_stat2trans = PENetwork_60_io_to_pes_14_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_190_io_data_1_in_valid = PENetwork_30_io_to_pes_14_in_valid; // @[pe.scala 264:34]
  assign PE_190_io_data_1_in_bits = PENetwork_30_io_to_pes_14_in_bits; // @[pe.scala 264:34]
  assign PE_190_io_data_0_in_valid = PENetwork_14_io_to_pes_8_in_valid; // @[pe.scala 264:34]
  assign PE_190_io_data_0_in_bits = PENetwork_14_io_to_pes_8_in_bits; // @[pe.scala 264:34]
  assign PE_191_clock = clock;
  assign PE_191_reset = reset;
  assign PE_191_io_data_2_sig_stat2trans = PENetwork_60_io_to_pes_15_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_191_io_data_1_in_valid = PENetwork_30_io_to_pes_15_in_valid; // @[pe.scala 264:34]
  assign PE_191_io_data_1_in_bits = PENetwork_30_io_to_pes_15_in_bits; // @[pe.scala 264:34]
  assign PE_191_io_data_0_in_valid = PENetwork_15_io_to_pes_8_in_valid; // @[pe.scala 264:34]
  assign PE_191_io_data_0_in_bits = PENetwork_15_io_to_pes_8_in_bits; // @[pe.scala 264:34]
  assign PE_192_clock = clock;
  assign PE_192_reset = reset;
  assign PE_192_io_data_2_sig_stat2trans = PENetwork_60_io_to_pes_16_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_192_io_data_1_in_valid = PENetwork_30_io_to_pes_16_in_valid; // @[pe.scala 264:34]
  assign PE_192_io_data_1_in_bits = PENetwork_30_io_to_pes_16_in_bits; // @[pe.scala 264:34]
  assign PE_192_io_data_0_in_valid = PENetwork_16_io_to_pes_8_in_valid; // @[pe.scala 264:34]
  assign PE_192_io_data_0_in_bits = PENetwork_16_io_to_pes_8_in_bits; // @[pe.scala 264:34]
  assign PE_193_clock = clock;
  assign PE_193_reset = reset;
  assign PE_193_io_data_2_sig_stat2trans = PENetwork_60_io_to_pes_17_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_193_io_data_1_in_valid = PENetwork_30_io_to_pes_17_in_valid; // @[pe.scala 264:34]
  assign PE_193_io_data_1_in_bits = PENetwork_30_io_to_pes_17_in_bits; // @[pe.scala 264:34]
  assign PE_193_io_data_0_in_valid = PENetwork_17_io_to_pes_8_in_valid; // @[pe.scala 264:34]
  assign PE_193_io_data_0_in_bits = PENetwork_17_io_to_pes_8_in_bits; // @[pe.scala 264:34]
  assign PE_194_clock = clock;
  assign PE_194_reset = reset;
  assign PE_194_io_data_2_sig_stat2trans = PENetwork_60_io_to_pes_18_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_194_io_data_1_in_valid = PENetwork_30_io_to_pes_18_in_valid; // @[pe.scala 264:34]
  assign PE_194_io_data_1_in_bits = PENetwork_30_io_to_pes_18_in_bits; // @[pe.scala 264:34]
  assign PE_194_io_data_0_in_valid = PENetwork_18_io_to_pes_8_in_valid; // @[pe.scala 264:34]
  assign PE_194_io_data_0_in_bits = PENetwork_18_io_to_pes_8_in_bits; // @[pe.scala 264:34]
  assign PE_195_clock = clock;
  assign PE_195_reset = reset;
  assign PE_195_io_data_2_sig_stat2trans = PENetwork_60_io_to_pes_19_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_195_io_data_1_in_valid = PENetwork_30_io_to_pes_19_in_valid; // @[pe.scala 264:34]
  assign PE_195_io_data_1_in_bits = PENetwork_30_io_to_pes_19_in_bits; // @[pe.scala 264:34]
  assign PE_195_io_data_0_in_valid = PENetwork_19_io_to_pes_8_in_valid; // @[pe.scala 264:34]
  assign PE_195_io_data_0_in_bits = PENetwork_19_io_to_pes_8_in_bits; // @[pe.scala 264:34]
  assign PE_196_clock = clock;
  assign PE_196_reset = reset;
  assign PE_196_io_data_2_sig_stat2trans = PENetwork_60_io_to_pes_20_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_196_io_data_1_in_valid = PENetwork_30_io_to_pes_20_in_valid; // @[pe.scala 264:34]
  assign PE_196_io_data_1_in_bits = PENetwork_30_io_to_pes_20_in_bits; // @[pe.scala 264:34]
  assign PE_196_io_data_0_in_valid = PENetwork_20_io_to_pes_8_in_valid; // @[pe.scala 264:34]
  assign PE_196_io_data_0_in_bits = PENetwork_20_io_to_pes_8_in_bits; // @[pe.scala 264:34]
  assign PE_197_clock = clock;
  assign PE_197_reset = reset;
  assign PE_197_io_data_2_sig_stat2trans = PENetwork_60_io_to_pes_21_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_197_io_data_1_in_valid = PENetwork_30_io_to_pes_21_in_valid; // @[pe.scala 264:34]
  assign PE_197_io_data_1_in_bits = PENetwork_30_io_to_pes_21_in_bits; // @[pe.scala 264:34]
  assign PE_197_io_data_0_in_valid = PENetwork_21_io_to_pes_8_in_valid; // @[pe.scala 264:34]
  assign PE_197_io_data_0_in_bits = PENetwork_21_io_to_pes_8_in_bits; // @[pe.scala 264:34]
  assign PE_198_clock = clock;
  assign PE_198_reset = reset;
  assign PE_198_io_data_2_sig_stat2trans = PENetwork_61_io_to_pes_0_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_198_io_data_1_in_valid = PENetwork_31_io_to_pes_0_in_valid; // @[pe.scala 264:34]
  assign PE_198_io_data_1_in_bits = PENetwork_31_io_to_pes_0_in_bits; // @[pe.scala 264:34]
  assign PE_198_io_data_0_in_valid = PENetwork_io_to_pes_9_in_valid; // @[pe.scala 264:34]
  assign PE_198_io_data_0_in_bits = PENetwork_io_to_pes_9_in_bits; // @[pe.scala 264:34]
  assign PE_199_clock = clock;
  assign PE_199_reset = reset;
  assign PE_199_io_data_2_sig_stat2trans = PENetwork_61_io_to_pes_1_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_199_io_data_1_in_valid = PENetwork_31_io_to_pes_1_in_valid; // @[pe.scala 264:34]
  assign PE_199_io_data_1_in_bits = PENetwork_31_io_to_pes_1_in_bits; // @[pe.scala 264:34]
  assign PE_199_io_data_0_in_valid = PENetwork_1_io_to_pes_9_in_valid; // @[pe.scala 264:34]
  assign PE_199_io_data_0_in_bits = PENetwork_1_io_to_pes_9_in_bits; // @[pe.scala 264:34]
  assign PE_200_clock = clock;
  assign PE_200_reset = reset;
  assign PE_200_io_data_2_sig_stat2trans = PENetwork_61_io_to_pes_2_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_200_io_data_1_in_valid = PENetwork_31_io_to_pes_2_in_valid; // @[pe.scala 264:34]
  assign PE_200_io_data_1_in_bits = PENetwork_31_io_to_pes_2_in_bits; // @[pe.scala 264:34]
  assign PE_200_io_data_0_in_valid = PENetwork_2_io_to_pes_9_in_valid; // @[pe.scala 264:34]
  assign PE_200_io_data_0_in_bits = PENetwork_2_io_to_pes_9_in_bits; // @[pe.scala 264:34]
  assign PE_201_clock = clock;
  assign PE_201_reset = reset;
  assign PE_201_io_data_2_sig_stat2trans = PENetwork_61_io_to_pes_3_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_201_io_data_1_in_valid = PENetwork_31_io_to_pes_3_in_valid; // @[pe.scala 264:34]
  assign PE_201_io_data_1_in_bits = PENetwork_31_io_to_pes_3_in_bits; // @[pe.scala 264:34]
  assign PE_201_io_data_0_in_valid = PENetwork_3_io_to_pes_9_in_valid; // @[pe.scala 264:34]
  assign PE_201_io_data_0_in_bits = PENetwork_3_io_to_pes_9_in_bits; // @[pe.scala 264:34]
  assign PE_202_clock = clock;
  assign PE_202_reset = reset;
  assign PE_202_io_data_2_sig_stat2trans = PENetwork_61_io_to_pes_4_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_202_io_data_1_in_valid = PENetwork_31_io_to_pes_4_in_valid; // @[pe.scala 264:34]
  assign PE_202_io_data_1_in_bits = PENetwork_31_io_to_pes_4_in_bits; // @[pe.scala 264:34]
  assign PE_202_io_data_0_in_valid = PENetwork_4_io_to_pes_9_in_valid; // @[pe.scala 264:34]
  assign PE_202_io_data_0_in_bits = PENetwork_4_io_to_pes_9_in_bits; // @[pe.scala 264:34]
  assign PE_203_clock = clock;
  assign PE_203_reset = reset;
  assign PE_203_io_data_2_sig_stat2trans = PENetwork_61_io_to_pes_5_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_203_io_data_1_in_valid = PENetwork_31_io_to_pes_5_in_valid; // @[pe.scala 264:34]
  assign PE_203_io_data_1_in_bits = PENetwork_31_io_to_pes_5_in_bits; // @[pe.scala 264:34]
  assign PE_203_io_data_0_in_valid = PENetwork_5_io_to_pes_9_in_valid; // @[pe.scala 264:34]
  assign PE_203_io_data_0_in_bits = PENetwork_5_io_to_pes_9_in_bits; // @[pe.scala 264:34]
  assign PE_204_clock = clock;
  assign PE_204_reset = reset;
  assign PE_204_io_data_2_sig_stat2trans = PENetwork_61_io_to_pes_6_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_204_io_data_1_in_valid = PENetwork_31_io_to_pes_6_in_valid; // @[pe.scala 264:34]
  assign PE_204_io_data_1_in_bits = PENetwork_31_io_to_pes_6_in_bits; // @[pe.scala 264:34]
  assign PE_204_io_data_0_in_valid = PENetwork_6_io_to_pes_9_in_valid; // @[pe.scala 264:34]
  assign PE_204_io_data_0_in_bits = PENetwork_6_io_to_pes_9_in_bits; // @[pe.scala 264:34]
  assign PE_205_clock = clock;
  assign PE_205_reset = reset;
  assign PE_205_io_data_2_sig_stat2trans = PENetwork_61_io_to_pes_7_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_205_io_data_1_in_valid = PENetwork_31_io_to_pes_7_in_valid; // @[pe.scala 264:34]
  assign PE_205_io_data_1_in_bits = PENetwork_31_io_to_pes_7_in_bits; // @[pe.scala 264:34]
  assign PE_205_io_data_0_in_valid = PENetwork_7_io_to_pes_9_in_valid; // @[pe.scala 264:34]
  assign PE_205_io_data_0_in_bits = PENetwork_7_io_to_pes_9_in_bits; // @[pe.scala 264:34]
  assign PE_206_clock = clock;
  assign PE_206_reset = reset;
  assign PE_206_io_data_2_sig_stat2trans = PENetwork_61_io_to_pes_8_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_206_io_data_1_in_valid = PENetwork_31_io_to_pes_8_in_valid; // @[pe.scala 264:34]
  assign PE_206_io_data_1_in_bits = PENetwork_31_io_to_pes_8_in_bits; // @[pe.scala 264:34]
  assign PE_206_io_data_0_in_valid = PENetwork_8_io_to_pes_9_in_valid; // @[pe.scala 264:34]
  assign PE_206_io_data_0_in_bits = PENetwork_8_io_to_pes_9_in_bits; // @[pe.scala 264:34]
  assign PE_207_clock = clock;
  assign PE_207_reset = reset;
  assign PE_207_io_data_2_sig_stat2trans = PENetwork_61_io_to_pes_9_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_207_io_data_1_in_valid = PENetwork_31_io_to_pes_9_in_valid; // @[pe.scala 264:34]
  assign PE_207_io_data_1_in_bits = PENetwork_31_io_to_pes_9_in_bits; // @[pe.scala 264:34]
  assign PE_207_io_data_0_in_valid = PENetwork_9_io_to_pes_9_in_valid; // @[pe.scala 264:34]
  assign PE_207_io_data_0_in_bits = PENetwork_9_io_to_pes_9_in_bits; // @[pe.scala 264:34]
  assign PE_208_clock = clock;
  assign PE_208_reset = reset;
  assign PE_208_io_data_2_sig_stat2trans = PENetwork_61_io_to_pes_10_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_208_io_data_1_in_valid = PENetwork_31_io_to_pes_10_in_valid; // @[pe.scala 264:34]
  assign PE_208_io_data_1_in_bits = PENetwork_31_io_to_pes_10_in_bits; // @[pe.scala 264:34]
  assign PE_208_io_data_0_in_valid = PENetwork_10_io_to_pes_9_in_valid; // @[pe.scala 264:34]
  assign PE_208_io_data_0_in_bits = PENetwork_10_io_to_pes_9_in_bits; // @[pe.scala 264:34]
  assign PE_209_clock = clock;
  assign PE_209_reset = reset;
  assign PE_209_io_data_2_sig_stat2trans = PENetwork_61_io_to_pes_11_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_209_io_data_1_in_valid = PENetwork_31_io_to_pes_11_in_valid; // @[pe.scala 264:34]
  assign PE_209_io_data_1_in_bits = PENetwork_31_io_to_pes_11_in_bits; // @[pe.scala 264:34]
  assign PE_209_io_data_0_in_valid = PENetwork_11_io_to_pes_9_in_valid; // @[pe.scala 264:34]
  assign PE_209_io_data_0_in_bits = PENetwork_11_io_to_pes_9_in_bits; // @[pe.scala 264:34]
  assign PE_210_clock = clock;
  assign PE_210_reset = reset;
  assign PE_210_io_data_2_sig_stat2trans = PENetwork_61_io_to_pes_12_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_210_io_data_1_in_valid = PENetwork_31_io_to_pes_12_in_valid; // @[pe.scala 264:34]
  assign PE_210_io_data_1_in_bits = PENetwork_31_io_to_pes_12_in_bits; // @[pe.scala 264:34]
  assign PE_210_io_data_0_in_valid = PENetwork_12_io_to_pes_9_in_valid; // @[pe.scala 264:34]
  assign PE_210_io_data_0_in_bits = PENetwork_12_io_to_pes_9_in_bits; // @[pe.scala 264:34]
  assign PE_211_clock = clock;
  assign PE_211_reset = reset;
  assign PE_211_io_data_2_sig_stat2trans = PENetwork_61_io_to_pes_13_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_211_io_data_1_in_valid = PENetwork_31_io_to_pes_13_in_valid; // @[pe.scala 264:34]
  assign PE_211_io_data_1_in_bits = PENetwork_31_io_to_pes_13_in_bits; // @[pe.scala 264:34]
  assign PE_211_io_data_0_in_valid = PENetwork_13_io_to_pes_9_in_valid; // @[pe.scala 264:34]
  assign PE_211_io_data_0_in_bits = PENetwork_13_io_to_pes_9_in_bits; // @[pe.scala 264:34]
  assign PE_212_clock = clock;
  assign PE_212_reset = reset;
  assign PE_212_io_data_2_sig_stat2trans = PENetwork_61_io_to_pes_14_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_212_io_data_1_in_valid = PENetwork_31_io_to_pes_14_in_valid; // @[pe.scala 264:34]
  assign PE_212_io_data_1_in_bits = PENetwork_31_io_to_pes_14_in_bits; // @[pe.scala 264:34]
  assign PE_212_io_data_0_in_valid = PENetwork_14_io_to_pes_9_in_valid; // @[pe.scala 264:34]
  assign PE_212_io_data_0_in_bits = PENetwork_14_io_to_pes_9_in_bits; // @[pe.scala 264:34]
  assign PE_213_clock = clock;
  assign PE_213_reset = reset;
  assign PE_213_io_data_2_sig_stat2trans = PENetwork_61_io_to_pes_15_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_213_io_data_1_in_valid = PENetwork_31_io_to_pes_15_in_valid; // @[pe.scala 264:34]
  assign PE_213_io_data_1_in_bits = PENetwork_31_io_to_pes_15_in_bits; // @[pe.scala 264:34]
  assign PE_213_io_data_0_in_valid = PENetwork_15_io_to_pes_9_in_valid; // @[pe.scala 264:34]
  assign PE_213_io_data_0_in_bits = PENetwork_15_io_to_pes_9_in_bits; // @[pe.scala 264:34]
  assign PE_214_clock = clock;
  assign PE_214_reset = reset;
  assign PE_214_io_data_2_sig_stat2trans = PENetwork_61_io_to_pes_16_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_214_io_data_1_in_valid = PENetwork_31_io_to_pes_16_in_valid; // @[pe.scala 264:34]
  assign PE_214_io_data_1_in_bits = PENetwork_31_io_to_pes_16_in_bits; // @[pe.scala 264:34]
  assign PE_214_io_data_0_in_valid = PENetwork_16_io_to_pes_9_in_valid; // @[pe.scala 264:34]
  assign PE_214_io_data_0_in_bits = PENetwork_16_io_to_pes_9_in_bits; // @[pe.scala 264:34]
  assign PE_215_clock = clock;
  assign PE_215_reset = reset;
  assign PE_215_io_data_2_sig_stat2trans = PENetwork_61_io_to_pes_17_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_215_io_data_1_in_valid = PENetwork_31_io_to_pes_17_in_valid; // @[pe.scala 264:34]
  assign PE_215_io_data_1_in_bits = PENetwork_31_io_to_pes_17_in_bits; // @[pe.scala 264:34]
  assign PE_215_io_data_0_in_valid = PENetwork_17_io_to_pes_9_in_valid; // @[pe.scala 264:34]
  assign PE_215_io_data_0_in_bits = PENetwork_17_io_to_pes_9_in_bits; // @[pe.scala 264:34]
  assign PE_216_clock = clock;
  assign PE_216_reset = reset;
  assign PE_216_io_data_2_sig_stat2trans = PENetwork_61_io_to_pes_18_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_216_io_data_1_in_valid = PENetwork_31_io_to_pes_18_in_valid; // @[pe.scala 264:34]
  assign PE_216_io_data_1_in_bits = PENetwork_31_io_to_pes_18_in_bits; // @[pe.scala 264:34]
  assign PE_216_io_data_0_in_valid = PENetwork_18_io_to_pes_9_in_valid; // @[pe.scala 264:34]
  assign PE_216_io_data_0_in_bits = PENetwork_18_io_to_pes_9_in_bits; // @[pe.scala 264:34]
  assign PE_217_clock = clock;
  assign PE_217_reset = reset;
  assign PE_217_io_data_2_sig_stat2trans = PENetwork_61_io_to_pes_19_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_217_io_data_1_in_valid = PENetwork_31_io_to_pes_19_in_valid; // @[pe.scala 264:34]
  assign PE_217_io_data_1_in_bits = PENetwork_31_io_to_pes_19_in_bits; // @[pe.scala 264:34]
  assign PE_217_io_data_0_in_valid = PENetwork_19_io_to_pes_9_in_valid; // @[pe.scala 264:34]
  assign PE_217_io_data_0_in_bits = PENetwork_19_io_to_pes_9_in_bits; // @[pe.scala 264:34]
  assign PE_218_clock = clock;
  assign PE_218_reset = reset;
  assign PE_218_io_data_2_sig_stat2trans = PENetwork_61_io_to_pes_20_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_218_io_data_1_in_valid = PENetwork_31_io_to_pes_20_in_valid; // @[pe.scala 264:34]
  assign PE_218_io_data_1_in_bits = PENetwork_31_io_to_pes_20_in_bits; // @[pe.scala 264:34]
  assign PE_218_io_data_0_in_valid = PENetwork_20_io_to_pes_9_in_valid; // @[pe.scala 264:34]
  assign PE_218_io_data_0_in_bits = PENetwork_20_io_to_pes_9_in_bits; // @[pe.scala 264:34]
  assign PE_219_clock = clock;
  assign PE_219_reset = reset;
  assign PE_219_io_data_2_sig_stat2trans = PENetwork_61_io_to_pes_21_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_219_io_data_1_in_valid = PENetwork_31_io_to_pes_21_in_valid; // @[pe.scala 264:34]
  assign PE_219_io_data_1_in_bits = PENetwork_31_io_to_pes_21_in_bits; // @[pe.scala 264:34]
  assign PE_219_io_data_0_in_valid = PENetwork_21_io_to_pes_9_in_valid; // @[pe.scala 264:34]
  assign PE_219_io_data_0_in_bits = PENetwork_21_io_to_pes_9_in_bits; // @[pe.scala 264:34]
  assign PE_220_clock = clock;
  assign PE_220_reset = reset;
  assign PE_220_io_data_2_sig_stat2trans = PENetwork_62_io_to_pes_0_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_220_io_data_1_in_valid = PENetwork_32_io_to_pes_0_in_valid; // @[pe.scala 264:34]
  assign PE_220_io_data_1_in_bits = PENetwork_32_io_to_pes_0_in_bits; // @[pe.scala 264:34]
  assign PE_220_io_data_0_in_valid = PENetwork_io_to_pes_10_in_valid; // @[pe.scala 264:34]
  assign PE_220_io_data_0_in_bits = PENetwork_io_to_pes_10_in_bits; // @[pe.scala 264:34]
  assign PE_221_clock = clock;
  assign PE_221_reset = reset;
  assign PE_221_io_data_2_sig_stat2trans = PENetwork_62_io_to_pes_1_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_221_io_data_1_in_valid = PENetwork_32_io_to_pes_1_in_valid; // @[pe.scala 264:34]
  assign PE_221_io_data_1_in_bits = PENetwork_32_io_to_pes_1_in_bits; // @[pe.scala 264:34]
  assign PE_221_io_data_0_in_valid = PENetwork_1_io_to_pes_10_in_valid; // @[pe.scala 264:34]
  assign PE_221_io_data_0_in_bits = PENetwork_1_io_to_pes_10_in_bits; // @[pe.scala 264:34]
  assign PE_222_clock = clock;
  assign PE_222_reset = reset;
  assign PE_222_io_data_2_sig_stat2trans = PENetwork_62_io_to_pes_2_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_222_io_data_1_in_valid = PENetwork_32_io_to_pes_2_in_valid; // @[pe.scala 264:34]
  assign PE_222_io_data_1_in_bits = PENetwork_32_io_to_pes_2_in_bits; // @[pe.scala 264:34]
  assign PE_222_io_data_0_in_valid = PENetwork_2_io_to_pes_10_in_valid; // @[pe.scala 264:34]
  assign PE_222_io_data_0_in_bits = PENetwork_2_io_to_pes_10_in_bits; // @[pe.scala 264:34]
  assign PE_223_clock = clock;
  assign PE_223_reset = reset;
  assign PE_223_io_data_2_sig_stat2trans = PENetwork_62_io_to_pes_3_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_223_io_data_1_in_valid = PENetwork_32_io_to_pes_3_in_valid; // @[pe.scala 264:34]
  assign PE_223_io_data_1_in_bits = PENetwork_32_io_to_pes_3_in_bits; // @[pe.scala 264:34]
  assign PE_223_io_data_0_in_valid = PENetwork_3_io_to_pes_10_in_valid; // @[pe.scala 264:34]
  assign PE_223_io_data_0_in_bits = PENetwork_3_io_to_pes_10_in_bits; // @[pe.scala 264:34]
  assign PE_224_clock = clock;
  assign PE_224_reset = reset;
  assign PE_224_io_data_2_sig_stat2trans = PENetwork_62_io_to_pes_4_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_224_io_data_1_in_valid = PENetwork_32_io_to_pes_4_in_valid; // @[pe.scala 264:34]
  assign PE_224_io_data_1_in_bits = PENetwork_32_io_to_pes_4_in_bits; // @[pe.scala 264:34]
  assign PE_224_io_data_0_in_valid = PENetwork_4_io_to_pes_10_in_valid; // @[pe.scala 264:34]
  assign PE_224_io_data_0_in_bits = PENetwork_4_io_to_pes_10_in_bits; // @[pe.scala 264:34]
  assign PE_225_clock = clock;
  assign PE_225_reset = reset;
  assign PE_225_io_data_2_sig_stat2trans = PENetwork_62_io_to_pes_5_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_225_io_data_1_in_valid = PENetwork_32_io_to_pes_5_in_valid; // @[pe.scala 264:34]
  assign PE_225_io_data_1_in_bits = PENetwork_32_io_to_pes_5_in_bits; // @[pe.scala 264:34]
  assign PE_225_io_data_0_in_valid = PENetwork_5_io_to_pes_10_in_valid; // @[pe.scala 264:34]
  assign PE_225_io_data_0_in_bits = PENetwork_5_io_to_pes_10_in_bits; // @[pe.scala 264:34]
  assign PE_226_clock = clock;
  assign PE_226_reset = reset;
  assign PE_226_io_data_2_sig_stat2trans = PENetwork_62_io_to_pes_6_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_226_io_data_1_in_valid = PENetwork_32_io_to_pes_6_in_valid; // @[pe.scala 264:34]
  assign PE_226_io_data_1_in_bits = PENetwork_32_io_to_pes_6_in_bits; // @[pe.scala 264:34]
  assign PE_226_io_data_0_in_valid = PENetwork_6_io_to_pes_10_in_valid; // @[pe.scala 264:34]
  assign PE_226_io_data_0_in_bits = PENetwork_6_io_to_pes_10_in_bits; // @[pe.scala 264:34]
  assign PE_227_clock = clock;
  assign PE_227_reset = reset;
  assign PE_227_io_data_2_sig_stat2trans = PENetwork_62_io_to_pes_7_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_227_io_data_1_in_valid = PENetwork_32_io_to_pes_7_in_valid; // @[pe.scala 264:34]
  assign PE_227_io_data_1_in_bits = PENetwork_32_io_to_pes_7_in_bits; // @[pe.scala 264:34]
  assign PE_227_io_data_0_in_valid = PENetwork_7_io_to_pes_10_in_valid; // @[pe.scala 264:34]
  assign PE_227_io_data_0_in_bits = PENetwork_7_io_to_pes_10_in_bits; // @[pe.scala 264:34]
  assign PE_228_clock = clock;
  assign PE_228_reset = reset;
  assign PE_228_io_data_2_sig_stat2trans = PENetwork_62_io_to_pes_8_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_228_io_data_1_in_valid = PENetwork_32_io_to_pes_8_in_valid; // @[pe.scala 264:34]
  assign PE_228_io_data_1_in_bits = PENetwork_32_io_to_pes_8_in_bits; // @[pe.scala 264:34]
  assign PE_228_io_data_0_in_valid = PENetwork_8_io_to_pes_10_in_valid; // @[pe.scala 264:34]
  assign PE_228_io_data_0_in_bits = PENetwork_8_io_to_pes_10_in_bits; // @[pe.scala 264:34]
  assign PE_229_clock = clock;
  assign PE_229_reset = reset;
  assign PE_229_io_data_2_sig_stat2trans = PENetwork_62_io_to_pes_9_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_229_io_data_1_in_valid = PENetwork_32_io_to_pes_9_in_valid; // @[pe.scala 264:34]
  assign PE_229_io_data_1_in_bits = PENetwork_32_io_to_pes_9_in_bits; // @[pe.scala 264:34]
  assign PE_229_io_data_0_in_valid = PENetwork_9_io_to_pes_10_in_valid; // @[pe.scala 264:34]
  assign PE_229_io_data_0_in_bits = PENetwork_9_io_to_pes_10_in_bits; // @[pe.scala 264:34]
  assign PE_230_clock = clock;
  assign PE_230_reset = reset;
  assign PE_230_io_data_2_sig_stat2trans = PENetwork_62_io_to_pes_10_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_230_io_data_1_in_valid = PENetwork_32_io_to_pes_10_in_valid; // @[pe.scala 264:34]
  assign PE_230_io_data_1_in_bits = PENetwork_32_io_to_pes_10_in_bits; // @[pe.scala 264:34]
  assign PE_230_io_data_0_in_valid = PENetwork_10_io_to_pes_10_in_valid; // @[pe.scala 264:34]
  assign PE_230_io_data_0_in_bits = PENetwork_10_io_to_pes_10_in_bits; // @[pe.scala 264:34]
  assign PE_231_clock = clock;
  assign PE_231_reset = reset;
  assign PE_231_io_data_2_sig_stat2trans = PENetwork_62_io_to_pes_11_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_231_io_data_1_in_valid = PENetwork_32_io_to_pes_11_in_valid; // @[pe.scala 264:34]
  assign PE_231_io_data_1_in_bits = PENetwork_32_io_to_pes_11_in_bits; // @[pe.scala 264:34]
  assign PE_231_io_data_0_in_valid = PENetwork_11_io_to_pes_10_in_valid; // @[pe.scala 264:34]
  assign PE_231_io_data_0_in_bits = PENetwork_11_io_to_pes_10_in_bits; // @[pe.scala 264:34]
  assign PE_232_clock = clock;
  assign PE_232_reset = reset;
  assign PE_232_io_data_2_sig_stat2trans = PENetwork_62_io_to_pes_12_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_232_io_data_1_in_valid = PENetwork_32_io_to_pes_12_in_valid; // @[pe.scala 264:34]
  assign PE_232_io_data_1_in_bits = PENetwork_32_io_to_pes_12_in_bits; // @[pe.scala 264:34]
  assign PE_232_io_data_0_in_valid = PENetwork_12_io_to_pes_10_in_valid; // @[pe.scala 264:34]
  assign PE_232_io_data_0_in_bits = PENetwork_12_io_to_pes_10_in_bits; // @[pe.scala 264:34]
  assign PE_233_clock = clock;
  assign PE_233_reset = reset;
  assign PE_233_io_data_2_sig_stat2trans = PENetwork_62_io_to_pes_13_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_233_io_data_1_in_valid = PENetwork_32_io_to_pes_13_in_valid; // @[pe.scala 264:34]
  assign PE_233_io_data_1_in_bits = PENetwork_32_io_to_pes_13_in_bits; // @[pe.scala 264:34]
  assign PE_233_io_data_0_in_valid = PENetwork_13_io_to_pes_10_in_valid; // @[pe.scala 264:34]
  assign PE_233_io_data_0_in_bits = PENetwork_13_io_to_pes_10_in_bits; // @[pe.scala 264:34]
  assign PE_234_clock = clock;
  assign PE_234_reset = reset;
  assign PE_234_io_data_2_sig_stat2trans = PENetwork_62_io_to_pes_14_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_234_io_data_1_in_valid = PENetwork_32_io_to_pes_14_in_valid; // @[pe.scala 264:34]
  assign PE_234_io_data_1_in_bits = PENetwork_32_io_to_pes_14_in_bits; // @[pe.scala 264:34]
  assign PE_234_io_data_0_in_valid = PENetwork_14_io_to_pes_10_in_valid; // @[pe.scala 264:34]
  assign PE_234_io_data_0_in_bits = PENetwork_14_io_to_pes_10_in_bits; // @[pe.scala 264:34]
  assign PE_235_clock = clock;
  assign PE_235_reset = reset;
  assign PE_235_io_data_2_sig_stat2trans = PENetwork_62_io_to_pes_15_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_235_io_data_1_in_valid = PENetwork_32_io_to_pes_15_in_valid; // @[pe.scala 264:34]
  assign PE_235_io_data_1_in_bits = PENetwork_32_io_to_pes_15_in_bits; // @[pe.scala 264:34]
  assign PE_235_io_data_0_in_valid = PENetwork_15_io_to_pes_10_in_valid; // @[pe.scala 264:34]
  assign PE_235_io_data_0_in_bits = PENetwork_15_io_to_pes_10_in_bits; // @[pe.scala 264:34]
  assign PE_236_clock = clock;
  assign PE_236_reset = reset;
  assign PE_236_io_data_2_sig_stat2trans = PENetwork_62_io_to_pes_16_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_236_io_data_1_in_valid = PENetwork_32_io_to_pes_16_in_valid; // @[pe.scala 264:34]
  assign PE_236_io_data_1_in_bits = PENetwork_32_io_to_pes_16_in_bits; // @[pe.scala 264:34]
  assign PE_236_io_data_0_in_valid = PENetwork_16_io_to_pes_10_in_valid; // @[pe.scala 264:34]
  assign PE_236_io_data_0_in_bits = PENetwork_16_io_to_pes_10_in_bits; // @[pe.scala 264:34]
  assign PE_237_clock = clock;
  assign PE_237_reset = reset;
  assign PE_237_io_data_2_sig_stat2trans = PENetwork_62_io_to_pes_17_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_237_io_data_1_in_valid = PENetwork_32_io_to_pes_17_in_valid; // @[pe.scala 264:34]
  assign PE_237_io_data_1_in_bits = PENetwork_32_io_to_pes_17_in_bits; // @[pe.scala 264:34]
  assign PE_237_io_data_0_in_valid = PENetwork_17_io_to_pes_10_in_valid; // @[pe.scala 264:34]
  assign PE_237_io_data_0_in_bits = PENetwork_17_io_to_pes_10_in_bits; // @[pe.scala 264:34]
  assign PE_238_clock = clock;
  assign PE_238_reset = reset;
  assign PE_238_io_data_2_sig_stat2trans = PENetwork_62_io_to_pes_18_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_238_io_data_1_in_valid = PENetwork_32_io_to_pes_18_in_valid; // @[pe.scala 264:34]
  assign PE_238_io_data_1_in_bits = PENetwork_32_io_to_pes_18_in_bits; // @[pe.scala 264:34]
  assign PE_238_io_data_0_in_valid = PENetwork_18_io_to_pes_10_in_valid; // @[pe.scala 264:34]
  assign PE_238_io_data_0_in_bits = PENetwork_18_io_to_pes_10_in_bits; // @[pe.scala 264:34]
  assign PE_239_clock = clock;
  assign PE_239_reset = reset;
  assign PE_239_io_data_2_sig_stat2trans = PENetwork_62_io_to_pes_19_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_239_io_data_1_in_valid = PENetwork_32_io_to_pes_19_in_valid; // @[pe.scala 264:34]
  assign PE_239_io_data_1_in_bits = PENetwork_32_io_to_pes_19_in_bits; // @[pe.scala 264:34]
  assign PE_239_io_data_0_in_valid = PENetwork_19_io_to_pes_10_in_valid; // @[pe.scala 264:34]
  assign PE_239_io_data_0_in_bits = PENetwork_19_io_to_pes_10_in_bits; // @[pe.scala 264:34]
  assign PE_240_clock = clock;
  assign PE_240_reset = reset;
  assign PE_240_io_data_2_sig_stat2trans = PENetwork_62_io_to_pes_20_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_240_io_data_1_in_valid = PENetwork_32_io_to_pes_20_in_valid; // @[pe.scala 264:34]
  assign PE_240_io_data_1_in_bits = PENetwork_32_io_to_pes_20_in_bits; // @[pe.scala 264:34]
  assign PE_240_io_data_0_in_valid = PENetwork_20_io_to_pes_10_in_valid; // @[pe.scala 264:34]
  assign PE_240_io_data_0_in_bits = PENetwork_20_io_to_pes_10_in_bits; // @[pe.scala 264:34]
  assign PE_241_clock = clock;
  assign PE_241_reset = reset;
  assign PE_241_io_data_2_sig_stat2trans = PENetwork_62_io_to_pes_21_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_241_io_data_1_in_valid = PENetwork_32_io_to_pes_21_in_valid; // @[pe.scala 264:34]
  assign PE_241_io_data_1_in_bits = PENetwork_32_io_to_pes_21_in_bits; // @[pe.scala 264:34]
  assign PE_241_io_data_0_in_valid = PENetwork_21_io_to_pes_10_in_valid; // @[pe.scala 264:34]
  assign PE_241_io_data_0_in_bits = PENetwork_21_io_to_pes_10_in_bits; // @[pe.scala 264:34]
  assign PE_242_clock = clock;
  assign PE_242_reset = reset;
  assign PE_242_io_data_2_sig_stat2trans = PENetwork_63_io_to_pes_0_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_242_io_data_1_in_valid = PENetwork_33_io_to_pes_0_in_valid; // @[pe.scala 264:34]
  assign PE_242_io_data_1_in_bits = PENetwork_33_io_to_pes_0_in_bits; // @[pe.scala 264:34]
  assign PE_242_io_data_0_in_valid = PENetwork_io_to_pes_11_in_valid; // @[pe.scala 264:34]
  assign PE_242_io_data_0_in_bits = PENetwork_io_to_pes_11_in_bits; // @[pe.scala 264:34]
  assign PE_243_clock = clock;
  assign PE_243_reset = reset;
  assign PE_243_io_data_2_sig_stat2trans = PENetwork_63_io_to_pes_1_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_243_io_data_1_in_valid = PENetwork_33_io_to_pes_1_in_valid; // @[pe.scala 264:34]
  assign PE_243_io_data_1_in_bits = PENetwork_33_io_to_pes_1_in_bits; // @[pe.scala 264:34]
  assign PE_243_io_data_0_in_valid = PENetwork_1_io_to_pes_11_in_valid; // @[pe.scala 264:34]
  assign PE_243_io_data_0_in_bits = PENetwork_1_io_to_pes_11_in_bits; // @[pe.scala 264:34]
  assign PE_244_clock = clock;
  assign PE_244_reset = reset;
  assign PE_244_io_data_2_sig_stat2trans = PENetwork_63_io_to_pes_2_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_244_io_data_1_in_valid = PENetwork_33_io_to_pes_2_in_valid; // @[pe.scala 264:34]
  assign PE_244_io_data_1_in_bits = PENetwork_33_io_to_pes_2_in_bits; // @[pe.scala 264:34]
  assign PE_244_io_data_0_in_valid = PENetwork_2_io_to_pes_11_in_valid; // @[pe.scala 264:34]
  assign PE_244_io_data_0_in_bits = PENetwork_2_io_to_pes_11_in_bits; // @[pe.scala 264:34]
  assign PE_245_clock = clock;
  assign PE_245_reset = reset;
  assign PE_245_io_data_2_sig_stat2trans = PENetwork_63_io_to_pes_3_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_245_io_data_1_in_valid = PENetwork_33_io_to_pes_3_in_valid; // @[pe.scala 264:34]
  assign PE_245_io_data_1_in_bits = PENetwork_33_io_to_pes_3_in_bits; // @[pe.scala 264:34]
  assign PE_245_io_data_0_in_valid = PENetwork_3_io_to_pes_11_in_valid; // @[pe.scala 264:34]
  assign PE_245_io_data_0_in_bits = PENetwork_3_io_to_pes_11_in_bits; // @[pe.scala 264:34]
  assign PE_246_clock = clock;
  assign PE_246_reset = reset;
  assign PE_246_io_data_2_sig_stat2trans = PENetwork_63_io_to_pes_4_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_246_io_data_1_in_valid = PENetwork_33_io_to_pes_4_in_valid; // @[pe.scala 264:34]
  assign PE_246_io_data_1_in_bits = PENetwork_33_io_to_pes_4_in_bits; // @[pe.scala 264:34]
  assign PE_246_io_data_0_in_valid = PENetwork_4_io_to_pes_11_in_valid; // @[pe.scala 264:34]
  assign PE_246_io_data_0_in_bits = PENetwork_4_io_to_pes_11_in_bits; // @[pe.scala 264:34]
  assign PE_247_clock = clock;
  assign PE_247_reset = reset;
  assign PE_247_io_data_2_sig_stat2trans = PENetwork_63_io_to_pes_5_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_247_io_data_1_in_valid = PENetwork_33_io_to_pes_5_in_valid; // @[pe.scala 264:34]
  assign PE_247_io_data_1_in_bits = PENetwork_33_io_to_pes_5_in_bits; // @[pe.scala 264:34]
  assign PE_247_io_data_0_in_valid = PENetwork_5_io_to_pes_11_in_valid; // @[pe.scala 264:34]
  assign PE_247_io_data_0_in_bits = PENetwork_5_io_to_pes_11_in_bits; // @[pe.scala 264:34]
  assign PE_248_clock = clock;
  assign PE_248_reset = reset;
  assign PE_248_io_data_2_sig_stat2trans = PENetwork_63_io_to_pes_6_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_248_io_data_1_in_valid = PENetwork_33_io_to_pes_6_in_valid; // @[pe.scala 264:34]
  assign PE_248_io_data_1_in_bits = PENetwork_33_io_to_pes_6_in_bits; // @[pe.scala 264:34]
  assign PE_248_io_data_0_in_valid = PENetwork_6_io_to_pes_11_in_valid; // @[pe.scala 264:34]
  assign PE_248_io_data_0_in_bits = PENetwork_6_io_to_pes_11_in_bits; // @[pe.scala 264:34]
  assign PE_249_clock = clock;
  assign PE_249_reset = reset;
  assign PE_249_io_data_2_sig_stat2trans = PENetwork_63_io_to_pes_7_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_249_io_data_1_in_valid = PENetwork_33_io_to_pes_7_in_valid; // @[pe.scala 264:34]
  assign PE_249_io_data_1_in_bits = PENetwork_33_io_to_pes_7_in_bits; // @[pe.scala 264:34]
  assign PE_249_io_data_0_in_valid = PENetwork_7_io_to_pes_11_in_valid; // @[pe.scala 264:34]
  assign PE_249_io_data_0_in_bits = PENetwork_7_io_to_pes_11_in_bits; // @[pe.scala 264:34]
  assign PE_250_clock = clock;
  assign PE_250_reset = reset;
  assign PE_250_io_data_2_sig_stat2trans = PENetwork_63_io_to_pes_8_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_250_io_data_1_in_valid = PENetwork_33_io_to_pes_8_in_valid; // @[pe.scala 264:34]
  assign PE_250_io_data_1_in_bits = PENetwork_33_io_to_pes_8_in_bits; // @[pe.scala 264:34]
  assign PE_250_io_data_0_in_valid = PENetwork_8_io_to_pes_11_in_valid; // @[pe.scala 264:34]
  assign PE_250_io_data_0_in_bits = PENetwork_8_io_to_pes_11_in_bits; // @[pe.scala 264:34]
  assign PE_251_clock = clock;
  assign PE_251_reset = reset;
  assign PE_251_io_data_2_sig_stat2trans = PENetwork_63_io_to_pes_9_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_251_io_data_1_in_valid = PENetwork_33_io_to_pes_9_in_valid; // @[pe.scala 264:34]
  assign PE_251_io_data_1_in_bits = PENetwork_33_io_to_pes_9_in_bits; // @[pe.scala 264:34]
  assign PE_251_io_data_0_in_valid = PENetwork_9_io_to_pes_11_in_valid; // @[pe.scala 264:34]
  assign PE_251_io_data_0_in_bits = PENetwork_9_io_to_pes_11_in_bits; // @[pe.scala 264:34]
  assign PE_252_clock = clock;
  assign PE_252_reset = reset;
  assign PE_252_io_data_2_sig_stat2trans = PENetwork_63_io_to_pes_10_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_252_io_data_1_in_valid = PENetwork_33_io_to_pes_10_in_valid; // @[pe.scala 264:34]
  assign PE_252_io_data_1_in_bits = PENetwork_33_io_to_pes_10_in_bits; // @[pe.scala 264:34]
  assign PE_252_io_data_0_in_valid = PENetwork_10_io_to_pes_11_in_valid; // @[pe.scala 264:34]
  assign PE_252_io_data_0_in_bits = PENetwork_10_io_to_pes_11_in_bits; // @[pe.scala 264:34]
  assign PE_253_clock = clock;
  assign PE_253_reset = reset;
  assign PE_253_io_data_2_sig_stat2trans = PENetwork_63_io_to_pes_11_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_253_io_data_1_in_valid = PENetwork_33_io_to_pes_11_in_valid; // @[pe.scala 264:34]
  assign PE_253_io_data_1_in_bits = PENetwork_33_io_to_pes_11_in_bits; // @[pe.scala 264:34]
  assign PE_253_io_data_0_in_valid = PENetwork_11_io_to_pes_11_in_valid; // @[pe.scala 264:34]
  assign PE_253_io_data_0_in_bits = PENetwork_11_io_to_pes_11_in_bits; // @[pe.scala 264:34]
  assign PE_254_clock = clock;
  assign PE_254_reset = reset;
  assign PE_254_io_data_2_sig_stat2trans = PENetwork_63_io_to_pes_12_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_254_io_data_1_in_valid = PENetwork_33_io_to_pes_12_in_valid; // @[pe.scala 264:34]
  assign PE_254_io_data_1_in_bits = PENetwork_33_io_to_pes_12_in_bits; // @[pe.scala 264:34]
  assign PE_254_io_data_0_in_valid = PENetwork_12_io_to_pes_11_in_valid; // @[pe.scala 264:34]
  assign PE_254_io_data_0_in_bits = PENetwork_12_io_to_pes_11_in_bits; // @[pe.scala 264:34]
  assign PE_255_clock = clock;
  assign PE_255_reset = reset;
  assign PE_255_io_data_2_sig_stat2trans = PENetwork_63_io_to_pes_13_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_255_io_data_1_in_valid = PENetwork_33_io_to_pes_13_in_valid; // @[pe.scala 264:34]
  assign PE_255_io_data_1_in_bits = PENetwork_33_io_to_pes_13_in_bits; // @[pe.scala 264:34]
  assign PE_255_io_data_0_in_valid = PENetwork_13_io_to_pes_11_in_valid; // @[pe.scala 264:34]
  assign PE_255_io_data_0_in_bits = PENetwork_13_io_to_pes_11_in_bits; // @[pe.scala 264:34]
  assign PE_256_clock = clock;
  assign PE_256_reset = reset;
  assign PE_256_io_data_2_sig_stat2trans = PENetwork_63_io_to_pes_14_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_256_io_data_1_in_valid = PENetwork_33_io_to_pes_14_in_valid; // @[pe.scala 264:34]
  assign PE_256_io_data_1_in_bits = PENetwork_33_io_to_pes_14_in_bits; // @[pe.scala 264:34]
  assign PE_256_io_data_0_in_valid = PENetwork_14_io_to_pes_11_in_valid; // @[pe.scala 264:34]
  assign PE_256_io_data_0_in_bits = PENetwork_14_io_to_pes_11_in_bits; // @[pe.scala 264:34]
  assign PE_257_clock = clock;
  assign PE_257_reset = reset;
  assign PE_257_io_data_2_sig_stat2trans = PENetwork_63_io_to_pes_15_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_257_io_data_1_in_valid = PENetwork_33_io_to_pes_15_in_valid; // @[pe.scala 264:34]
  assign PE_257_io_data_1_in_bits = PENetwork_33_io_to_pes_15_in_bits; // @[pe.scala 264:34]
  assign PE_257_io_data_0_in_valid = PENetwork_15_io_to_pes_11_in_valid; // @[pe.scala 264:34]
  assign PE_257_io_data_0_in_bits = PENetwork_15_io_to_pes_11_in_bits; // @[pe.scala 264:34]
  assign PE_258_clock = clock;
  assign PE_258_reset = reset;
  assign PE_258_io_data_2_sig_stat2trans = PENetwork_63_io_to_pes_16_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_258_io_data_1_in_valid = PENetwork_33_io_to_pes_16_in_valid; // @[pe.scala 264:34]
  assign PE_258_io_data_1_in_bits = PENetwork_33_io_to_pes_16_in_bits; // @[pe.scala 264:34]
  assign PE_258_io_data_0_in_valid = PENetwork_16_io_to_pes_11_in_valid; // @[pe.scala 264:34]
  assign PE_258_io_data_0_in_bits = PENetwork_16_io_to_pes_11_in_bits; // @[pe.scala 264:34]
  assign PE_259_clock = clock;
  assign PE_259_reset = reset;
  assign PE_259_io_data_2_sig_stat2trans = PENetwork_63_io_to_pes_17_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_259_io_data_1_in_valid = PENetwork_33_io_to_pes_17_in_valid; // @[pe.scala 264:34]
  assign PE_259_io_data_1_in_bits = PENetwork_33_io_to_pes_17_in_bits; // @[pe.scala 264:34]
  assign PE_259_io_data_0_in_valid = PENetwork_17_io_to_pes_11_in_valid; // @[pe.scala 264:34]
  assign PE_259_io_data_0_in_bits = PENetwork_17_io_to_pes_11_in_bits; // @[pe.scala 264:34]
  assign PE_260_clock = clock;
  assign PE_260_reset = reset;
  assign PE_260_io_data_2_sig_stat2trans = PENetwork_63_io_to_pes_18_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_260_io_data_1_in_valid = PENetwork_33_io_to_pes_18_in_valid; // @[pe.scala 264:34]
  assign PE_260_io_data_1_in_bits = PENetwork_33_io_to_pes_18_in_bits; // @[pe.scala 264:34]
  assign PE_260_io_data_0_in_valid = PENetwork_18_io_to_pes_11_in_valid; // @[pe.scala 264:34]
  assign PE_260_io_data_0_in_bits = PENetwork_18_io_to_pes_11_in_bits; // @[pe.scala 264:34]
  assign PE_261_clock = clock;
  assign PE_261_reset = reset;
  assign PE_261_io_data_2_sig_stat2trans = PENetwork_63_io_to_pes_19_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_261_io_data_1_in_valid = PENetwork_33_io_to_pes_19_in_valid; // @[pe.scala 264:34]
  assign PE_261_io_data_1_in_bits = PENetwork_33_io_to_pes_19_in_bits; // @[pe.scala 264:34]
  assign PE_261_io_data_0_in_valid = PENetwork_19_io_to_pes_11_in_valid; // @[pe.scala 264:34]
  assign PE_261_io_data_0_in_bits = PENetwork_19_io_to_pes_11_in_bits; // @[pe.scala 264:34]
  assign PE_262_clock = clock;
  assign PE_262_reset = reset;
  assign PE_262_io_data_2_sig_stat2trans = PENetwork_63_io_to_pes_20_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_262_io_data_1_in_valid = PENetwork_33_io_to_pes_20_in_valid; // @[pe.scala 264:34]
  assign PE_262_io_data_1_in_bits = PENetwork_33_io_to_pes_20_in_bits; // @[pe.scala 264:34]
  assign PE_262_io_data_0_in_valid = PENetwork_20_io_to_pes_11_in_valid; // @[pe.scala 264:34]
  assign PE_262_io_data_0_in_bits = PENetwork_20_io_to_pes_11_in_bits; // @[pe.scala 264:34]
  assign PE_263_clock = clock;
  assign PE_263_reset = reset;
  assign PE_263_io_data_2_sig_stat2trans = PENetwork_63_io_to_pes_21_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_263_io_data_1_in_valid = PENetwork_33_io_to_pes_21_in_valid; // @[pe.scala 264:34]
  assign PE_263_io_data_1_in_bits = PENetwork_33_io_to_pes_21_in_bits; // @[pe.scala 264:34]
  assign PE_263_io_data_0_in_valid = PENetwork_21_io_to_pes_11_in_valid; // @[pe.scala 264:34]
  assign PE_263_io_data_0_in_bits = PENetwork_21_io_to_pes_11_in_bits; // @[pe.scala 264:34]
  assign PE_264_clock = clock;
  assign PE_264_reset = reset;
  assign PE_264_io_data_2_sig_stat2trans = PENetwork_64_io_to_pes_0_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_264_io_data_1_in_valid = PENetwork_34_io_to_pes_0_in_valid; // @[pe.scala 264:34]
  assign PE_264_io_data_1_in_bits = PENetwork_34_io_to_pes_0_in_bits; // @[pe.scala 264:34]
  assign PE_264_io_data_0_in_valid = PENetwork_io_to_pes_12_in_valid; // @[pe.scala 264:34]
  assign PE_264_io_data_0_in_bits = PENetwork_io_to_pes_12_in_bits; // @[pe.scala 264:34]
  assign PE_265_clock = clock;
  assign PE_265_reset = reset;
  assign PE_265_io_data_2_sig_stat2trans = PENetwork_64_io_to_pes_1_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_265_io_data_1_in_valid = PENetwork_34_io_to_pes_1_in_valid; // @[pe.scala 264:34]
  assign PE_265_io_data_1_in_bits = PENetwork_34_io_to_pes_1_in_bits; // @[pe.scala 264:34]
  assign PE_265_io_data_0_in_valid = PENetwork_1_io_to_pes_12_in_valid; // @[pe.scala 264:34]
  assign PE_265_io_data_0_in_bits = PENetwork_1_io_to_pes_12_in_bits; // @[pe.scala 264:34]
  assign PE_266_clock = clock;
  assign PE_266_reset = reset;
  assign PE_266_io_data_2_sig_stat2trans = PENetwork_64_io_to_pes_2_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_266_io_data_1_in_valid = PENetwork_34_io_to_pes_2_in_valid; // @[pe.scala 264:34]
  assign PE_266_io_data_1_in_bits = PENetwork_34_io_to_pes_2_in_bits; // @[pe.scala 264:34]
  assign PE_266_io_data_0_in_valid = PENetwork_2_io_to_pes_12_in_valid; // @[pe.scala 264:34]
  assign PE_266_io_data_0_in_bits = PENetwork_2_io_to_pes_12_in_bits; // @[pe.scala 264:34]
  assign PE_267_clock = clock;
  assign PE_267_reset = reset;
  assign PE_267_io_data_2_sig_stat2trans = PENetwork_64_io_to_pes_3_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_267_io_data_1_in_valid = PENetwork_34_io_to_pes_3_in_valid; // @[pe.scala 264:34]
  assign PE_267_io_data_1_in_bits = PENetwork_34_io_to_pes_3_in_bits; // @[pe.scala 264:34]
  assign PE_267_io_data_0_in_valid = PENetwork_3_io_to_pes_12_in_valid; // @[pe.scala 264:34]
  assign PE_267_io_data_0_in_bits = PENetwork_3_io_to_pes_12_in_bits; // @[pe.scala 264:34]
  assign PE_268_clock = clock;
  assign PE_268_reset = reset;
  assign PE_268_io_data_2_sig_stat2trans = PENetwork_64_io_to_pes_4_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_268_io_data_1_in_valid = PENetwork_34_io_to_pes_4_in_valid; // @[pe.scala 264:34]
  assign PE_268_io_data_1_in_bits = PENetwork_34_io_to_pes_4_in_bits; // @[pe.scala 264:34]
  assign PE_268_io_data_0_in_valid = PENetwork_4_io_to_pes_12_in_valid; // @[pe.scala 264:34]
  assign PE_268_io_data_0_in_bits = PENetwork_4_io_to_pes_12_in_bits; // @[pe.scala 264:34]
  assign PE_269_clock = clock;
  assign PE_269_reset = reset;
  assign PE_269_io_data_2_sig_stat2trans = PENetwork_64_io_to_pes_5_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_269_io_data_1_in_valid = PENetwork_34_io_to_pes_5_in_valid; // @[pe.scala 264:34]
  assign PE_269_io_data_1_in_bits = PENetwork_34_io_to_pes_5_in_bits; // @[pe.scala 264:34]
  assign PE_269_io_data_0_in_valid = PENetwork_5_io_to_pes_12_in_valid; // @[pe.scala 264:34]
  assign PE_269_io_data_0_in_bits = PENetwork_5_io_to_pes_12_in_bits; // @[pe.scala 264:34]
  assign PE_270_clock = clock;
  assign PE_270_reset = reset;
  assign PE_270_io_data_2_sig_stat2trans = PENetwork_64_io_to_pes_6_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_270_io_data_1_in_valid = PENetwork_34_io_to_pes_6_in_valid; // @[pe.scala 264:34]
  assign PE_270_io_data_1_in_bits = PENetwork_34_io_to_pes_6_in_bits; // @[pe.scala 264:34]
  assign PE_270_io_data_0_in_valid = PENetwork_6_io_to_pes_12_in_valid; // @[pe.scala 264:34]
  assign PE_270_io_data_0_in_bits = PENetwork_6_io_to_pes_12_in_bits; // @[pe.scala 264:34]
  assign PE_271_clock = clock;
  assign PE_271_reset = reset;
  assign PE_271_io_data_2_sig_stat2trans = PENetwork_64_io_to_pes_7_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_271_io_data_1_in_valid = PENetwork_34_io_to_pes_7_in_valid; // @[pe.scala 264:34]
  assign PE_271_io_data_1_in_bits = PENetwork_34_io_to_pes_7_in_bits; // @[pe.scala 264:34]
  assign PE_271_io_data_0_in_valid = PENetwork_7_io_to_pes_12_in_valid; // @[pe.scala 264:34]
  assign PE_271_io_data_0_in_bits = PENetwork_7_io_to_pes_12_in_bits; // @[pe.scala 264:34]
  assign PE_272_clock = clock;
  assign PE_272_reset = reset;
  assign PE_272_io_data_2_sig_stat2trans = PENetwork_64_io_to_pes_8_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_272_io_data_1_in_valid = PENetwork_34_io_to_pes_8_in_valid; // @[pe.scala 264:34]
  assign PE_272_io_data_1_in_bits = PENetwork_34_io_to_pes_8_in_bits; // @[pe.scala 264:34]
  assign PE_272_io_data_0_in_valid = PENetwork_8_io_to_pes_12_in_valid; // @[pe.scala 264:34]
  assign PE_272_io_data_0_in_bits = PENetwork_8_io_to_pes_12_in_bits; // @[pe.scala 264:34]
  assign PE_273_clock = clock;
  assign PE_273_reset = reset;
  assign PE_273_io_data_2_sig_stat2trans = PENetwork_64_io_to_pes_9_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_273_io_data_1_in_valid = PENetwork_34_io_to_pes_9_in_valid; // @[pe.scala 264:34]
  assign PE_273_io_data_1_in_bits = PENetwork_34_io_to_pes_9_in_bits; // @[pe.scala 264:34]
  assign PE_273_io_data_0_in_valid = PENetwork_9_io_to_pes_12_in_valid; // @[pe.scala 264:34]
  assign PE_273_io_data_0_in_bits = PENetwork_9_io_to_pes_12_in_bits; // @[pe.scala 264:34]
  assign PE_274_clock = clock;
  assign PE_274_reset = reset;
  assign PE_274_io_data_2_sig_stat2trans = PENetwork_64_io_to_pes_10_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_274_io_data_1_in_valid = PENetwork_34_io_to_pes_10_in_valid; // @[pe.scala 264:34]
  assign PE_274_io_data_1_in_bits = PENetwork_34_io_to_pes_10_in_bits; // @[pe.scala 264:34]
  assign PE_274_io_data_0_in_valid = PENetwork_10_io_to_pes_12_in_valid; // @[pe.scala 264:34]
  assign PE_274_io_data_0_in_bits = PENetwork_10_io_to_pes_12_in_bits; // @[pe.scala 264:34]
  assign PE_275_clock = clock;
  assign PE_275_reset = reset;
  assign PE_275_io_data_2_sig_stat2trans = PENetwork_64_io_to_pes_11_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_275_io_data_1_in_valid = PENetwork_34_io_to_pes_11_in_valid; // @[pe.scala 264:34]
  assign PE_275_io_data_1_in_bits = PENetwork_34_io_to_pes_11_in_bits; // @[pe.scala 264:34]
  assign PE_275_io_data_0_in_valid = PENetwork_11_io_to_pes_12_in_valid; // @[pe.scala 264:34]
  assign PE_275_io_data_0_in_bits = PENetwork_11_io_to_pes_12_in_bits; // @[pe.scala 264:34]
  assign PE_276_clock = clock;
  assign PE_276_reset = reset;
  assign PE_276_io_data_2_sig_stat2trans = PENetwork_64_io_to_pes_12_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_276_io_data_1_in_valid = PENetwork_34_io_to_pes_12_in_valid; // @[pe.scala 264:34]
  assign PE_276_io_data_1_in_bits = PENetwork_34_io_to_pes_12_in_bits; // @[pe.scala 264:34]
  assign PE_276_io_data_0_in_valid = PENetwork_12_io_to_pes_12_in_valid; // @[pe.scala 264:34]
  assign PE_276_io_data_0_in_bits = PENetwork_12_io_to_pes_12_in_bits; // @[pe.scala 264:34]
  assign PE_277_clock = clock;
  assign PE_277_reset = reset;
  assign PE_277_io_data_2_sig_stat2trans = PENetwork_64_io_to_pes_13_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_277_io_data_1_in_valid = PENetwork_34_io_to_pes_13_in_valid; // @[pe.scala 264:34]
  assign PE_277_io_data_1_in_bits = PENetwork_34_io_to_pes_13_in_bits; // @[pe.scala 264:34]
  assign PE_277_io_data_0_in_valid = PENetwork_13_io_to_pes_12_in_valid; // @[pe.scala 264:34]
  assign PE_277_io_data_0_in_bits = PENetwork_13_io_to_pes_12_in_bits; // @[pe.scala 264:34]
  assign PE_278_clock = clock;
  assign PE_278_reset = reset;
  assign PE_278_io_data_2_sig_stat2trans = PENetwork_64_io_to_pes_14_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_278_io_data_1_in_valid = PENetwork_34_io_to_pes_14_in_valid; // @[pe.scala 264:34]
  assign PE_278_io_data_1_in_bits = PENetwork_34_io_to_pes_14_in_bits; // @[pe.scala 264:34]
  assign PE_278_io_data_0_in_valid = PENetwork_14_io_to_pes_12_in_valid; // @[pe.scala 264:34]
  assign PE_278_io_data_0_in_bits = PENetwork_14_io_to_pes_12_in_bits; // @[pe.scala 264:34]
  assign PE_279_clock = clock;
  assign PE_279_reset = reset;
  assign PE_279_io_data_2_sig_stat2trans = PENetwork_64_io_to_pes_15_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_279_io_data_1_in_valid = PENetwork_34_io_to_pes_15_in_valid; // @[pe.scala 264:34]
  assign PE_279_io_data_1_in_bits = PENetwork_34_io_to_pes_15_in_bits; // @[pe.scala 264:34]
  assign PE_279_io_data_0_in_valid = PENetwork_15_io_to_pes_12_in_valid; // @[pe.scala 264:34]
  assign PE_279_io_data_0_in_bits = PENetwork_15_io_to_pes_12_in_bits; // @[pe.scala 264:34]
  assign PE_280_clock = clock;
  assign PE_280_reset = reset;
  assign PE_280_io_data_2_sig_stat2trans = PENetwork_64_io_to_pes_16_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_280_io_data_1_in_valid = PENetwork_34_io_to_pes_16_in_valid; // @[pe.scala 264:34]
  assign PE_280_io_data_1_in_bits = PENetwork_34_io_to_pes_16_in_bits; // @[pe.scala 264:34]
  assign PE_280_io_data_0_in_valid = PENetwork_16_io_to_pes_12_in_valid; // @[pe.scala 264:34]
  assign PE_280_io_data_0_in_bits = PENetwork_16_io_to_pes_12_in_bits; // @[pe.scala 264:34]
  assign PE_281_clock = clock;
  assign PE_281_reset = reset;
  assign PE_281_io_data_2_sig_stat2trans = PENetwork_64_io_to_pes_17_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_281_io_data_1_in_valid = PENetwork_34_io_to_pes_17_in_valid; // @[pe.scala 264:34]
  assign PE_281_io_data_1_in_bits = PENetwork_34_io_to_pes_17_in_bits; // @[pe.scala 264:34]
  assign PE_281_io_data_0_in_valid = PENetwork_17_io_to_pes_12_in_valid; // @[pe.scala 264:34]
  assign PE_281_io_data_0_in_bits = PENetwork_17_io_to_pes_12_in_bits; // @[pe.scala 264:34]
  assign PE_282_clock = clock;
  assign PE_282_reset = reset;
  assign PE_282_io_data_2_sig_stat2trans = PENetwork_64_io_to_pes_18_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_282_io_data_1_in_valid = PENetwork_34_io_to_pes_18_in_valid; // @[pe.scala 264:34]
  assign PE_282_io_data_1_in_bits = PENetwork_34_io_to_pes_18_in_bits; // @[pe.scala 264:34]
  assign PE_282_io_data_0_in_valid = PENetwork_18_io_to_pes_12_in_valid; // @[pe.scala 264:34]
  assign PE_282_io_data_0_in_bits = PENetwork_18_io_to_pes_12_in_bits; // @[pe.scala 264:34]
  assign PE_283_clock = clock;
  assign PE_283_reset = reset;
  assign PE_283_io_data_2_sig_stat2trans = PENetwork_64_io_to_pes_19_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_283_io_data_1_in_valid = PENetwork_34_io_to_pes_19_in_valid; // @[pe.scala 264:34]
  assign PE_283_io_data_1_in_bits = PENetwork_34_io_to_pes_19_in_bits; // @[pe.scala 264:34]
  assign PE_283_io_data_0_in_valid = PENetwork_19_io_to_pes_12_in_valid; // @[pe.scala 264:34]
  assign PE_283_io_data_0_in_bits = PENetwork_19_io_to_pes_12_in_bits; // @[pe.scala 264:34]
  assign PE_284_clock = clock;
  assign PE_284_reset = reset;
  assign PE_284_io_data_2_sig_stat2trans = PENetwork_64_io_to_pes_20_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_284_io_data_1_in_valid = PENetwork_34_io_to_pes_20_in_valid; // @[pe.scala 264:34]
  assign PE_284_io_data_1_in_bits = PENetwork_34_io_to_pes_20_in_bits; // @[pe.scala 264:34]
  assign PE_284_io_data_0_in_valid = PENetwork_20_io_to_pes_12_in_valid; // @[pe.scala 264:34]
  assign PE_284_io_data_0_in_bits = PENetwork_20_io_to_pes_12_in_bits; // @[pe.scala 264:34]
  assign PE_285_clock = clock;
  assign PE_285_reset = reset;
  assign PE_285_io_data_2_sig_stat2trans = PENetwork_64_io_to_pes_21_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_285_io_data_1_in_valid = PENetwork_34_io_to_pes_21_in_valid; // @[pe.scala 264:34]
  assign PE_285_io_data_1_in_bits = PENetwork_34_io_to_pes_21_in_bits; // @[pe.scala 264:34]
  assign PE_285_io_data_0_in_valid = PENetwork_21_io_to_pes_12_in_valid; // @[pe.scala 264:34]
  assign PE_285_io_data_0_in_bits = PENetwork_21_io_to_pes_12_in_bits; // @[pe.scala 264:34]
  assign PE_286_clock = clock;
  assign PE_286_reset = reset;
  assign PE_286_io_data_2_sig_stat2trans = PENetwork_65_io_to_pes_0_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_286_io_data_1_in_valid = PENetwork_35_io_to_pes_0_in_valid; // @[pe.scala 264:34]
  assign PE_286_io_data_1_in_bits = PENetwork_35_io_to_pes_0_in_bits; // @[pe.scala 264:34]
  assign PE_286_io_data_0_in_valid = PENetwork_io_to_pes_13_in_valid; // @[pe.scala 264:34]
  assign PE_286_io_data_0_in_bits = PENetwork_io_to_pes_13_in_bits; // @[pe.scala 264:34]
  assign PE_287_clock = clock;
  assign PE_287_reset = reset;
  assign PE_287_io_data_2_sig_stat2trans = PENetwork_65_io_to_pes_1_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_287_io_data_1_in_valid = PENetwork_35_io_to_pes_1_in_valid; // @[pe.scala 264:34]
  assign PE_287_io_data_1_in_bits = PENetwork_35_io_to_pes_1_in_bits; // @[pe.scala 264:34]
  assign PE_287_io_data_0_in_valid = PENetwork_1_io_to_pes_13_in_valid; // @[pe.scala 264:34]
  assign PE_287_io_data_0_in_bits = PENetwork_1_io_to_pes_13_in_bits; // @[pe.scala 264:34]
  assign PE_288_clock = clock;
  assign PE_288_reset = reset;
  assign PE_288_io_data_2_sig_stat2trans = PENetwork_65_io_to_pes_2_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_288_io_data_1_in_valid = PENetwork_35_io_to_pes_2_in_valid; // @[pe.scala 264:34]
  assign PE_288_io_data_1_in_bits = PENetwork_35_io_to_pes_2_in_bits; // @[pe.scala 264:34]
  assign PE_288_io_data_0_in_valid = PENetwork_2_io_to_pes_13_in_valid; // @[pe.scala 264:34]
  assign PE_288_io_data_0_in_bits = PENetwork_2_io_to_pes_13_in_bits; // @[pe.scala 264:34]
  assign PE_289_clock = clock;
  assign PE_289_reset = reset;
  assign PE_289_io_data_2_sig_stat2trans = PENetwork_65_io_to_pes_3_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_289_io_data_1_in_valid = PENetwork_35_io_to_pes_3_in_valid; // @[pe.scala 264:34]
  assign PE_289_io_data_1_in_bits = PENetwork_35_io_to_pes_3_in_bits; // @[pe.scala 264:34]
  assign PE_289_io_data_0_in_valid = PENetwork_3_io_to_pes_13_in_valid; // @[pe.scala 264:34]
  assign PE_289_io_data_0_in_bits = PENetwork_3_io_to_pes_13_in_bits; // @[pe.scala 264:34]
  assign PE_290_clock = clock;
  assign PE_290_reset = reset;
  assign PE_290_io_data_2_sig_stat2trans = PENetwork_65_io_to_pes_4_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_290_io_data_1_in_valid = PENetwork_35_io_to_pes_4_in_valid; // @[pe.scala 264:34]
  assign PE_290_io_data_1_in_bits = PENetwork_35_io_to_pes_4_in_bits; // @[pe.scala 264:34]
  assign PE_290_io_data_0_in_valid = PENetwork_4_io_to_pes_13_in_valid; // @[pe.scala 264:34]
  assign PE_290_io_data_0_in_bits = PENetwork_4_io_to_pes_13_in_bits; // @[pe.scala 264:34]
  assign PE_291_clock = clock;
  assign PE_291_reset = reset;
  assign PE_291_io_data_2_sig_stat2trans = PENetwork_65_io_to_pes_5_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_291_io_data_1_in_valid = PENetwork_35_io_to_pes_5_in_valid; // @[pe.scala 264:34]
  assign PE_291_io_data_1_in_bits = PENetwork_35_io_to_pes_5_in_bits; // @[pe.scala 264:34]
  assign PE_291_io_data_0_in_valid = PENetwork_5_io_to_pes_13_in_valid; // @[pe.scala 264:34]
  assign PE_291_io_data_0_in_bits = PENetwork_5_io_to_pes_13_in_bits; // @[pe.scala 264:34]
  assign PE_292_clock = clock;
  assign PE_292_reset = reset;
  assign PE_292_io_data_2_sig_stat2trans = PENetwork_65_io_to_pes_6_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_292_io_data_1_in_valid = PENetwork_35_io_to_pes_6_in_valid; // @[pe.scala 264:34]
  assign PE_292_io_data_1_in_bits = PENetwork_35_io_to_pes_6_in_bits; // @[pe.scala 264:34]
  assign PE_292_io_data_0_in_valid = PENetwork_6_io_to_pes_13_in_valid; // @[pe.scala 264:34]
  assign PE_292_io_data_0_in_bits = PENetwork_6_io_to_pes_13_in_bits; // @[pe.scala 264:34]
  assign PE_293_clock = clock;
  assign PE_293_reset = reset;
  assign PE_293_io_data_2_sig_stat2trans = PENetwork_65_io_to_pes_7_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_293_io_data_1_in_valid = PENetwork_35_io_to_pes_7_in_valid; // @[pe.scala 264:34]
  assign PE_293_io_data_1_in_bits = PENetwork_35_io_to_pes_7_in_bits; // @[pe.scala 264:34]
  assign PE_293_io_data_0_in_valid = PENetwork_7_io_to_pes_13_in_valid; // @[pe.scala 264:34]
  assign PE_293_io_data_0_in_bits = PENetwork_7_io_to_pes_13_in_bits; // @[pe.scala 264:34]
  assign PE_294_clock = clock;
  assign PE_294_reset = reset;
  assign PE_294_io_data_2_sig_stat2trans = PENetwork_65_io_to_pes_8_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_294_io_data_1_in_valid = PENetwork_35_io_to_pes_8_in_valid; // @[pe.scala 264:34]
  assign PE_294_io_data_1_in_bits = PENetwork_35_io_to_pes_8_in_bits; // @[pe.scala 264:34]
  assign PE_294_io_data_0_in_valid = PENetwork_8_io_to_pes_13_in_valid; // @[pe.scala 264:34]
  assign PE_294_io_data_0_in_bits = PENetwork_8_io_to_pes_13_in_bits; // @[pe.scala 264:34]
  assign PE_295_clock = clock;
  assign PE_295_reset = reset;
  assign PE_295_io_data_2_sig_stat2trans = PENetwork_65_io_to_pes_9_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_295_io_data_1_in_valid = PENetwork_35_io_to_pes_9_in_valid; // @[pe.scala 264:34]
  assign PE_295_io_data_1_in_bits = PENetwork_35_io_to_pes_9_in_bits; // @[pe.scala 264:34]
  assign PE_295_io_data_0_in_valid = PENetwork_9_io_to_pes_13_in_valid; // @[pe.scala 264:34]
  assign PE_295_io_data_0_in_bits = PENetwork_9_io_to_pes_13_in_bits; // @[pe.scala 264:34]
  assign PE_296_clock = clock;
  assign PE_296_reset = reset;
  assign PE_296_io_data_2_sig_stat2trans = PENetwork_65_io_to_pes_10_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_296_io_data_1_in_valid = PENetwork_35_io_to_pes_10_in_valid; // @[pe.scala 264:34]
  assign PE_296_io_data_1_in_bits = PENetwork_35_io_to_pes_10_in_bits; // @[pe.scala 264:34]
  assign PE_296_io_data_0_in_valid = PENetwork_10_io_to_pes_13_in_valid; // @[pe.scala 264:34]
  assign PE_296_io_data_0_in_bits = PENetwork_10_io_to_pes_13_in_bits; // @[pe.scala 264:34]
  assign PE_297_clock = clock;
  assign PE_297_reset = reset;
  assign PE_297_io_data_2_sig_stat2trans = PENetwork_65_io_to_pes_11_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_297_io_data_1_in_valid = PENetwork_35_io_to_pes_11_in_valid; // @[pe.scala 264:34]
  assign PE_297_io_data_1_in_bits = PENetwork_35_io_to_pes_11_in_bits; // @[pe.scala 264:34]
  assign PE_297_io_data_0_in_valid = PENetwork_11_io_to_pes_13_in_valid; // @[pe.scala 264:34]
  assign PE_297_io_data_0_in_bits = PENetwork_11_io_to_pes_13_in_bits; // @[pe.scala 264:34]
  assign PE_298_clock = clock;
  assign PE_298_reset = reset;
  assign PE_298_io_data_2_sig_stat2trans = PENetwork_65_io_to_pes_12_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_298_io_data_1_in_valid = PENetwork_35_io_to_pes_12_in_valid; // @[pe.scala 264:34]
  assign PE_298_io_data_1_in_bits = PENetwork_35_io_to_pes_12_in_bits; // @[pe.scala 264:34]
  assign PE_298_io_data_0_in_valid = PENetwork_12_io_to_pes_13_in_valid; // @[pe.scala 264:34]
  assign PE_298_io_data_0_in_bits = PENetwork_12_io_to_pes_13_in_bits; // @[pe.scala 264:34]
  assign PE_299_clock = clock;
  assign PE_299_reset = reset;
  assign PE_299_io_data_2_sig_stat2trans = PENetwork_65_io_to_pes_13_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_299_io_data_1_in_valid = PENetwork_35_io_to_pes_13_in_valid; // @[pe.scala 264:34]
  assign PE_299_io_data_1_in_bits = PENetwork_35_io_to_pes_13_in_bits; // @[pe.scala 264:34]
  assign PE_299_io_data_0_in_valid = PENetwork_13_io_to_pes_13_in_valid; // @[pe.scala 264:34]
  assign PE_299_io_data_0_in_bits = PENetwork_13_io_to_pes_13_in_bits; // @[pe.scala 264:34]
  assign PE_300_clock = clock;
  assign PE_300_reset = reset;
  assign PE_300_io_data_2_sig_stat2trans = PENetwork_65_io_to_pes_14_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_300_io_data_1_in_valid = PENetwork_35_io_to_pes_14_in_valid; // @[pe.scala 264:34]
  assign PE_300_io_data_1_in_bits = PENetwork_35_io_to_pes_14_in_bits; // @[pe.scala 264:34]
  assign PE_300_io_data_0_in_valid = PENetwork_14_io_to_pes_13_in_valid; // @[pe.scala 264:34]
  assign PE_300_io_data_0_in_bits = PENetwork_14_io_to_pes_13_in_bits; // @[pe.scala 264:34]
  assign PE_301_clock = clock;
  assign PE_301_reset = reset;
  assign PE_301_io_data_2_sig_stat2trans = PENetwork_65_io_to_pes_15_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_301_io_data_1_in_valid = PENetwork_35_io_to_pes_15_in_valid; // @[pe.scala 264:34]
  assign PE_301_io_data_1_in_bits = PENetwork_35_io_to_pes_15_in_bits; // @[pe.scala 264:34]
  assign PE_301_io_data_0_in_valid = PENetwork_15_io_to_pes_13_in_valid; // @[pe.scala 264:34]
  assign PE_301_io_data_0_in_bits = PENetwork_15_io_to_pes_13_in_bits; // @[pe.scala 264:34]
  assign PE_302_clock = clock;
  assign PE_302_reset = reset;
  assign PE_302_io_data_2_sig_stat2trans = PENetwork_65_io_to_pes_16_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_302_io_data_1_in_valid = PENetwork_35_io_to_pes_16_in_valid; // @[pe.scala 264:34]
  assign PE_302_io_data_1_in_bits = PENetwork_35_io_to_pes_16_in_bits; // @[pe.scala 264:34]
  assign PE_302_io_data_0_in_valid = PENetwork_16_io_to_pes_13_in_valid; // @[pe.scala 264:34]
  assign PE_302_io_data_0_in_bits = PENetwork_16_io_to_pes_13_in_bits; // @[pe.scala 264:34]
  assign PE_303_clock = clock;
  assign PE_303_reset = reset;
  assign PE_303_io_data_2_sig_stat2trans = PENetwork_65_io_to_pes_17_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_303_io_data_1_in_valid = PENetwork_35_io_to_pes_17_in_valid; // @[pe.scala 264:34]
  assign PE_303_io_data_1_in_bits = PENetwork_35_io_to_pes_17_in_bits; // @[pe.scala 264:34]
  assign PE_303_io_data_0_in_valid = PENetwork_17_io_to_pes_13_in_valid; // @[pe.scala 264:34]
  assign PE_303_io_data_0_in_bits = PENetwork_17_io_to_pes_13_in_bits; // @[pe.scala 264:34]
  assign PE_304_clock = clock;
  assign PE_304_reset = reset;
  assign PE_304_io_data_2_sig_stat2trans = PENetwork_65_io_to_pes_18_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_304_io_data_1_in_valid = PENetwork_35_io_to_pes_18_in_valid; // @[pe.scala 264:34]
  assign PE_304_io_data_1_in_bits = PENetwork_35_io_to_pes_18_in_bits; // @[pe.scala 264:34]
  assign PE_304_io_data_0_in_valid = PENetwork_18_io_to_pes_13_in_valid; // @[pe.scala 264:34]
  assign PE_304_io_data_0_in_bits = PENetwork_18_io_to_pes_13_in_bits; // @[pe.scala 264:34]
  assign PE_305_clock = clock;
  assign PE_305_reset = reset;
  assign PE_305_io_data_2_sig_stat2trans = PENetwork_65_io_to_pes_19_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_305_io_data_1_in_valid = PENetwork_35_io_to_pes_19_in_valid; // @[pe.scala 264:34]
  assign PE_305_io_data_1_in_bits = PENetwork_35_io_to_pes_19_in_bits; // @[pe.scala 264:34]
  assign PE_305_io_data_0_in_valid = PENetwork_19_io_to_pes_13_in_valid; // @[pe.scala 264:34]
  assign PE_305_io_data_0_in_bits = PENetwork_19_io_to_pes_13_in_bits; // @[pe.scala 264:34]
  assign PE_306_clock = clock;
  assign PE_306_reset = reset;
  assign PE_306_io_data_2_sig_stat2trans = PENetwork_65_io_to_pes_20_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_306_io_data_1_in_valid = PENetwork_35_io_to_pes_20_in_valid; // @[pe.scala 264:34]
  assign PE_306_io_data_1_in_bits = PENetwork_35_io_to_pes_20_in_bits; // @[pe.scala 264:34]
  assign PE_306_io_data_0_in_valid = PENetwork_20_io_to_pes_13_in_valid; // @[pe.scala 264:34]
  assign PE_306_io_data_0_in_bits = PENetwork_20_io_to_pes_13_in_bits; // @[pe.scala 264:34]
  assign PE_307_clock = clock;
  assign PE_307_reset = reset;
  assign PE_307_io_data_2_sig_stat2trans = PENetwork_65_io_to_pes_21_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_307_io_data_1_in_valid = PENetwork_35_io_to_pes_21_in_valid; // @[pe.scala 264:34]
  assign PE_307_io_data_1_in_bits = PENetwork_35_io_to_pes_21_in_bits; // @[pe.scala 264:34]
  assign PE_307_io_data_0_in_valid = PENetwork_21_io_to_pes_13_in_valid; // @[pe.scala 264:34]
  assign PE_307_io_data_0_in_bits = PENetwork_21_io_to_pes_13_in_bits; // @[pe.scala 264:34]
  assign PE_308_clock = clock;
  assign PE_308_reset = reset;
  assign PE_308_io_data_2_sig_stat2trans = PENetwork_66_io_to_pes_0_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_308_io_data_1_in_valid = PENetwork_36_io_to_pes_0_in_valid; // @[pe.scala 264:34]
  assign PE_308_io_data_1_in_bits = PENetwork_36_io_to_pes_0_in_bits; // @[pe.scala 264:34]
  assign PE_308_io_data_0_in_valid = PENetwork_io_to_pes_14_in_valid; // @[pe.scala 264:34]
  assign PE_308_io_data_0_in_bits = PENetwork_io_to_pes_14_in_bits; // @[pe.scala 264:34]
  assign PE_309_clock = clock;
  assign PE_309_reset = reset;
  assign PE_309_io_data_2_sig_stat2trans = PENetwork_66_io_to_pes_1_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_309_io_data_1_in_valid = PENetwork_36_io_to_pes_1_in_valid; // @[pe.scala 264:34]
  assign PE_309_io_data_1_in_bits = PENetwork_36_io_to_pes_1_in_bits; // @[pe.scala 264:34]
  assign PE_309_io_data_0_in_valid = PENetwork_1_io_to_pes_14_in_valid; // @[pe.scala 264:34]
  assign PE_309_io_data_0_in_bits = PENetwork_1_io_to_pes_14_in_bits; // @[pe.scala 264:34]
  assign PE_310_clock = clock;
  assign PE_310_reset = reset;
  assign PE_310_io_data_2_sig_stat2trans = PENetwork_66_io_to_pes_2_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_310_io_data_1_in_valid = PENetwork_36_io_to_pes_2_in_valid; // @[pe.scala 264:34]
  assign PE_310_io_data_1_in_bits = PENetwork_36_io_to_pes_2_in_bits; // @[pe.scala 264:34]
  assign PE_310_io_data_0_in_valid = PENetwork_2_io_to_pes_14_in_valid; // @[pe.scala 264:34]
  assign PE_310_io_data_0_in_bits = PENetwork_2_io_to_pes_14_in_bits; // @[pe.scala 264:34]
  assign PE_311_clock = clock;
  assign PE_311_reset = reset;
  assign PE_311_io_data_2_sig_stat2trans = PENetwork_66_io_to_pes_3_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_311_io_data_1_in_valid = PENetwork_36_io_to_pes_3_in_valid; // @[pe.scala 264:34]
  assign PE_311_io_data_1_in_bits = PENetwork_36_io_to_pes_3_in_bits; // @[pe.scala 264:34]
  assign PE_311_io_data_0_in_valid = PENetwork_3_io_to_pes_14_in_valid; // @[pe.scala 264:34]
  assign PE_311_io_data_0_in_bits = PENetwork_3_io_to_pes_14_in_bits; // @[pe.scala 264:34]
  assign PE_312_clock = clock;
  assign PE_312_reset = reset;
  assign PE_312_io_data_2_sig_stat2trans = PENetwork_66_io_to_pes_4_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_312_io_data_1_in_valid = PENetwork_36_io_to_pes_4_in_valid; // @[pe.scala 264:34]
  assign PE_312_io_data_1_in_bits = PENetwork_36_io_to_pes_4_in_bits; // @[pe.scala 264:34]
  assign PE_312_io_data_0_in_valid = PENetwork_4_io_to_pes_14_in_valid; // @[pe.scala 264:34]
  assign PE_312_io_data_0_in_bits = PENetwork_4_io_to_pes_14_in_bits; // @[pe.scala 264:34]
  assign PE_313_clock = clock;
  assign PE_313_reset = reset;
  assign PE_313_io_data_2_sig_stat2trans = PENetwork_66_io_to_pes_5_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_313_io_data_1_in_valid = PENetwork_36_io_to_pes_5_in_valid; // @[pe.scala 264:34]
  assign PE_313_io_data_1_in_bits = PENetwork_36_io_to_pes_5_in_bits; // @[pe.scala 264:34]
  assign PE_313_io_data_0_in_valid = PENetwork_5_io_to_pes_14_in_valid; // @[pe.scala 264:34]
  assign PE_313_io_data_0_in_bits = PENetwork_5_io_to_pes_14_in_bits; // @[pe.scala 264:34]
  assign PE_314_clock = clock;
  assign PE_314_reset = reset;
  assign PE_314_io_data_2_sig_stat2trans = PENetwork_66_io_to_pes_6_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_314_io_data_1_in_valid = PENetwork_36_io_to_pes_6_in_valid; // @[pe.scala 264:34]
  assign PE_314_io_data_1_in_bits = PENetwork_36_io_to_pes_6_in_bits; // @[pe.scala 264:34]
  assign PE_314_io_data_0_in_valid = PENetwork_6_io_to_pes_14_in_valid; // @[pe.scala 264:34]
  assign PE_314_io_data_0_in_bits = PENetwork_6_io_to_pes_14_in_bits; // @[pe.scala 264:34]
  assign PE_315_clock = clock;
  assign PE_315_reset = reset;
  assign PE_315_io_data_2_sig_stat2trans = PENetwork_66_io_to_pes_7_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_315_io_data_1_in_valid = PENetwork_36_io_to_pes_7_in_valid; // @[pe.scala 264:34]
  assign PE_315_io_data_1_in_bits = PENetwork_36_io_to_pes_7_in_bits; // @[pe.scala 264:34]
  assign PE_315_io_data_0_in_valid = PENetwork_7_io_to_pes_14_in_valid; // @[pe.scala 264:34]
  assign PE_315_io_data_0_in_bits = PENetwork_7_io_to_pes_14_in_bits; // @[pe.scala 264:34]
  assign PE_316_clock = clock;
  assign PE_316_reset = reset;
  assign PE_316_io_data_2_sig_stat2trans = PENetwork_66_io_to_pes_8_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_316_io_data_1_in_valid = PENetwork_36_io_to_pes_8_in_valid; // @[pe.scala 264:34]
  assign PE_316_io_data_1_in_bits = PENetwork_36_io_to_pes_8_in_bits; // @[pe.scala 264:34]
  assign PE_316_io_data_0_in_valid = PENetwork_8_io_to_pes_14_in_valid; // @[pe.scala 264:34]
  assign PE_316_io_data_0_in_bits = PENetwork_8_io_to_pes_14_in_bits; // @[pe.scala 264:34]
  assign PE_317_clock = clock;
  assign PE_317_reset = reset;
  assign PE_317_io_data_2_sig_stat2trans = PENetwork_66_io_to_pes_9_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_317_io_data_1_in_valid = PENetwork_36_io_to_pes_9_in_valid; // @[pe.scala 264:34]
  assign PE_317_io_data_1_in_bits = PENetwork_36_io_to_pes_9_in_bits; // @[pe.scala 264:34]
  assign PE_317_io_data_0_in_valid = PENetwork_9_io_to_pes_14_in_valid; // @[pe.scala 264:34]
  assign PE_317_io_data_0_in_bits = PENetwork_9_io_to_pes_14_in_bits; // @[pe.scala 264:34]
  assign PE_318_clock = clock;
  assign PE_318_reset = reset;
  assign PE_318_io_data_2_sig_stat2trans = PENetwork_66_io_to_pes_10_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_318_io_data_1_in_valid = PENetwork_36_io_to_pes_10_in_valid; // @[pe.scala 264:34]
  assign PE_318_io_data_1_in_bits = PENetwork_36_io_to_pes_10_in_bits; // @[pe.scala 264:34]
  assign PE_318_io_data_0_in_valid = PENetwork_10_io_to_pes_14_in_valid; // @[pe.scala 264:34]
  assign PE_318_io_data_0_in_bits = PENetwork_10_io_to_pes_14_in_bits; // @[pe.scala 264:34]
  assign PE_319_clock = clock;
  assign PE_319_reset = reset;
  assign PE_319_io_data_2_sig_stat2trans = PENetwork_66_io_to_pes_11_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_319_io_data_1_in_valid = PENetwork_36_io_to_pes_11_in_valid; // @[pe.scala 264:34]
  assign PE_319_io_data_1_in_bits = PENetwork_36_io_to_pes_11_in_bits; // @[pe.scala 264:34]
  assign PE_319_io_data_0_in_valid = PENetwork_11_io_to_pes_14_in_valid; // @[pe.scala 264:34]
  assign PE_319_io_data_0_in_bits = PENetwork_11_io_to_pes_14_in_bits; // @[pe.scala 264:34]
  assign PE_320_clock = clock;
  assign PE_320_reset = reset;
  assign PE_320_io_data_2_sig_stat2trans = PENetwork_66_io_to_pes_12_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_320_io_data_1_in_valid = PENetwork_36_io_to_pes_12_in_valid; // @[pe.scala 264:34]
  assign PE_320_io_data_1_in_bits = PENetwork_36_io_to_pes_12_in_bits; // @[pe.scala 264:34]
  assign PE_320_io_data_0_in_valid = PENetwork_12_io_to_pes_14_in_valid; // @[pe.scala 264:34]
  assign PE_320_io_data_0_in_bits = PENetwork_12_io_to_pes_14_in_bits; // @[pe.scala 264:34]
  assign PE_321_clock = clock;
  assign PE_321_reset = reset;
  assign PE_321_io_data_2_sig_stat2trans = PENetwork_66_io_to_pes_13_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_321_io_data_1_in_valid = PENetwork_36_io_to_pes_13_in_valid; // @[pe.scala 264:34]
  assign PE_321_io_data_1_in_bits = PENetwork_36_io_to_pes_13_in_bits; // @[pe.scala 264:34]
  assign PE_321_io_data_0_in_valid = PENetwork_13_io_to_pes_14_in_valid; // @[pe.scala 264:34]
  assign PE_321_io_data_0_in_bits = PENetwork_13_io_to_pes_14_in_bits; // @[pe.scala 264:34]
  assign PE_322_clock = clock;
  assign PE_322_reset = reset;
  assign PE_322_io_data_2_sig_stat2trans = PENetwork_66_io_to_pes_14_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_322_io_data_1_in_valid = PENetwork_36_io_to_pes_14_in_valid; // @[pe.scala 264:34]
  assign PE_322_io_data_1_in_bits = PENetwork_36_io_to_pes_14_in_bits; // @[pe.scala 264:34]
  assign PE_322_io_data_0_in_valid = PENetwork_14_io_to_pes_14_in_valid; // @[pe.scala 264:34]
  assign PE_322_io_data_0_in_bits = PENetwork_14_io_to_pes_14_in_bits; // @[pe.scala 264:34]
  assign PE_323_clock = clock;
  assign PE_323_reset = reset;
  assign PE_323_io_data_2_sig_stat2trans = PENetwork_66_io_to_pes_15_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_323_io_data_1_in_valid = PENetwork_36_io_to_pes_15_in_valid; // @[pe.scala 264:34]
  assign PE_323_io_data_1_in_bits = PENetwork_36_io_to_pes_15_in_bits; // @[pe.scala 264:34]
  assign PE_323_io_data_0_in_valid = PENetwork_15_io_to_pes_14_in_valid; // @[pe.scala 264:34]
  assign PE_323_io_data_0_in_bits = PENetwork_15_io_to_pes_14_in_bits; // @[pe.scala 264:34]
  assign PE_324_clock = clock;
  assign PE_324_reset = reset;
  assign PE_324_io_data_2_sig_stat2trans = PENetwork_66_io_to_pes_16_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_324_io_data_1_in_valid = PENetwork_36_io_to_pes_16_in_valid; // @[pe.scala 264:34]
  assign PE_324_io_data_1_in_bits = PENetwork_36_io_to_pes_16_in_bits; // @[pe.scala 264:34]
  assign PE_324_io_data_0_in_valid = PENetwork_16_io_to_pes_14_in_valid; // @[pe.scala 264:34]
  assign PE_324_io_data_0_in_bits = PENetwork_16_io_to_pes_14_in_bits; // @[pe.scala 264:34]
  assign PE_325_clock = clock;
  assign PE_325_reset = reset;
  assign PE_325_io_data_2_sig_stat2trans = PENetwork_66_io_to_pes_17_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_325_io_data_1_in_valid = PENetwork_36_io_to_pes_17_in_valid; // @[pe.scala 264:34]
  assign PE_325_io_data_1_in_bits = PENetwork_36_io_to_pes_17_in_bits; // @[pe.scala 264:34]
  assign PE_325_io_data_0_in_valid = PENetwork_17_io_to_pes_14_in_valid; // @[pe.scala 264:34]
  assign PE_325_io_data_0_in_bits = PENetwork_17_io_to_pes_14_in_bits; // @[pe.scala 264:34]
  assign PE_326_clock = clock;
  assign PE_326_reset = reset;
  assign PE_326_io_data_2_sig_stat2trans = PENetwork_66_io_to_pes_18_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_326_io_data_1_in_valid = PENetwork_36_io_to_pes_18_in_valid; // @[pe.scala 264:34]
  assign PE_326_io_data_1_in_bits = PENetwork_36_io_to_pes_18_in_bits; // @[pe.scala 264:34]
  assign PE_326_io_data_0_in_valid = PENetwork_18_io_to_pes_14_in_valid; // @[pe.scala 264:34]
  assign PE_326_io_data_0_in_bits = PENetwork_18_io_to_pes_14_in_bits; // @[pe.scala 264:34]
  assign PE_327_clock = clock;
  assign PE_327_reset = reset;
  assign PE_327_io_data_2_sig_stat2trans = PENetwork_66_io_to_pes_19_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_327_io_data_1_in_valid = PENetwork_36_io_to_pes_19_in_valid; // @[pe.scala 264:34]
  assign PE_327_io_data_1_in_bits = PENetwork_36_io_to_pes_19_in_bits; // @[pe.scala 264:34]
  assign PE_327_io_data_0_in_valid = PENetwork_19_io_to_pes_14_in_valid; // @[pe.scala 264:34]
  assign PE_327_io_data_0_in_bits = PENetwork_19_io_to_pes_14_in_bits; // @[pe.scala 264:34]
  assign PE_328_clock = clock;
  assign PE_328_reset = reset;
  assign PE_328_io_data_2_sig_stat2trans = PENetwork_66_io_to_pes_20_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_328_io_data_1_in_valid = PENetwork_36_io_to_pes_20_in_valid; // @[pe.scala 264:34]
  assign PE_328_io_data_1_in_bits = PENetwork_36_io_to_pes_20_in_bits; // @[pe.scala 264:34]
  assign PE_328_io_data_0_in_valid = PENetwork_20_io_to_pes_14_in_valid; // @[pe.scala 264:34]
  assign PE_328_io_data_0_in_bits = PENetwork_20_io_to_pes_14_in_bits; // @[pe.scala 264:34]
  assign PE_329_clock = clock;
  assign PE_329_reset = reset;
  assign PE_329_io_data_2_sig_stat2trans = PENetwork_66_io_to_pes_21_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_329_io_data_1_in_valid = PENetwork_36_io_to_pes_21_in_valid; // @[pe.scala 264:34]
  assign PE_329_io_data_1_in_bits = PENetwork_36_io_to_pes_21_in_bits; // @[pe.scala 264:34]
  assign PE_329_io_data_0_in_valid = PENetwork_21_io_to_pes_14_in_valid; // @[pe.scala 264:34]
  assign PE_329_io_data_0_in_bits = PENetwork_21_io_to_pes_14_in_bits; // @[pe.scala 264:34]
  assign PE_330_clock = clock;
  assign PE_330_reset = reset;
  assign PE_330_io_data_2_sig_stat2trans = PENetwork_67_io_to_pes_0_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_330_io_data_1_in_valid = PENetwork_37_io_to_pes_0_in_valid; // @[pe.scala 264:34]
  assign PE_330_io_data_1_in_bits = PENetwork_37_io_to_pes_0_in_bits; // @[pe.scala 264:34]
  assign PE_330_io_data_0_in_valid = PENetwork_io_to_pes_15_in_valid; // @[pe.scala 264:34]
  assign PE_330_io_data_0_in_bits = PENetwork_io_to_pes_15_in_bits; // @[pe.scala 264:34]
  assign PE_331_clock = clock;
  assign PE_331_reset = reset;
  assign PE_331_io_data_2_sig_stat2trans = PENetwork_67_io_to_pes_1_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_331_io_data_1_in_valid = PENetwork_37_io_to_pes_1_in_valid; // @[pe.scala 264:34]
  assign PE_331_io_data_1_in_bits = PENetwork_37_io_to_pes_1_in_bits; // @[pe.scala 264:34]
  assign PE_331_io_data_0_in_valid = PENetwork_1_io_to_pes_15_in_valid; // @[pe.scala 264:34]
  assign PE_331_io_data_0_in_bits = PENetwork_1_io_to_pes_15_in_bits; // @[pe.scala 264:34]
  assign PE_332_clock = clock;
  assign PE_332_reset = reset;
  assign PE_332_io_data_2_sig_stat2trans = PENetwork_67_io_to_pes_2_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_332_io_data_1_in_valid = PENetwork_37_io_to_pes_2_in_valid; // @[pe.scala 264:34]
  assign PE_332_io_data_1_in_bits = PENetwork_37_io_to_pes_2_in_bits; // @[pe.scala 264:34]
  assign PE_332_io_data_0_in_valid = PENetwork_2_io_to_pes_15_in_valid; // @[pe.scala 264:34]
  assign PE_332_io_data_0_in_bits = PENetwork_2_io_to_pes_15_in_bits; // @[pe.scala 264:34]
  assign PE_333_clock = clock;
  assign PE_333_reset = reset;
  assign PE_333_io_data_2_sig_stat2trans = PENetwork_67_io_to_pes_3_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_333_io_data_1_in_valid = PENetwork_37_io_to_pes_3_in_valid; // @[pe.scala 264:34]
  assign PE_333_io_data_1_in_bits = PENetwork_37_io_to_pes_3_in_bits; // @[pe.scala 264:34]
  assign PE_333_io_data_0_in_valid = PENetwork_3_io_to_pes_15_in_valid; // @[pe.scala 264:34]
  assign PE_333_io_data_0_in_bits = PENetwork_3_io_to_pes_15_in_bits; // @[pe.scala 264:34]
  assign PE_334_clock = clock;
  assign PE_334_reset = reset;
  assign PE_334_io_data_2_sig_stat2trans = PENetwork_67_io_to_pes_4_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_334_io_data_1_in_valid = PENetwork_37_io_to_pes_4_in_valid; // @[pe.scala 264:34]
  assign PE_334_io_data_1_in_bits = PENetwork_37_io_to_pes_4_in_bits; // @[pe.scala 264:34]
  assign PE_334_io_data_0_in_valid = PENetwork_4_io_to_pes_15_in_valid; // @[pe.scala 264:34]
  assign PE_334_io_data_0_in_bits = PENetwork_4_io_to_pes_15_in_bits; // @[pe.scala 264:34]
  assign PE_335_clock = clock;
  assign PE_335_reset = reset;
  assign PE_335_io_data_2_sig_stat2trans = PENetwork_67_io_to_pes_5_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_335_io_data_1_in_valid = PENetwork_37_io_to_pes_5_in_valid; // @[pe.scala 264:34]
  assign PE_335_io_data_1_in_bits = PENetwork_37_io_to_pes_5_in_bits; // @[pe.scala 264:34]
  assign PE_335_io_data_0_in_valid = PENetwork_5_io_to_pes_15_in_valid; // @[pe.scala 264:34]
  assign PE_335_io_data_0_in_bits = PENetwork_5_io_to_pes_15_in_bits; // @[pe.scala 264:34]
  assign PE_336_clock = clock;
  assign PE_336_reset = reset;
  assign PE_336_io_data_2_sig_stat2trans = PENetwork_67_io_to_pes_6_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_336_io_data_1_in_valid = PENetwork_37_io_to_pes_6_in_valid; // @[pe.scala 264:34]
  assign PE_336_io_data_1_in_bits = PENetwork_37_io_to_pes_6_in_bits; // @[pe.scala 264:34]
  assign PE_336_io_data_0_in_valid = PENetwork_6_io_to_pes_15_in_valid; // @[pe.scala 264:34]
  assign PE_336_io_data_0_in_bits = PENetwork_6_io_to_pes_15_in_bits; // @[pe.scala 264:34]
  assign PE_337_clock = clock;
  assign PE_337_reset = reset;
  assign PE_337_io_data_2_sig_stat2trans = PENetwork_67_io_to_pes_7_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_337_io_data_1_in_valid = PENetwork_37_io_to_pes_7_in_valid; // @[pe.scala 264:34]
  assign PE_337_io_data_1_in_bits = PENetwork_37_io_to_pes_7_in_bits; // @[pe.scala 264:34]
  assign PE_337_io_data_0_in_valid = PENetwork_7_io_to_pes_15_in_valid; // @[pe.scala 264:34]
  assign PE_337_io_data_0_in_bits = PENetwork_7_io_to_pes_15_in_bits; // @[pe.scala 264:34]
  assign PE_338_clock = clock;
  assign PE_338_reset = reset;
  assign PE_338_io_data_2_sig_stat2trans = PENetwork_67_io_to_pes_8_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_338_io_data_1_in_valid = PENetwork_37_io_to_pes_8_in_valid; // @[pe.scala 264:34]
  assign PE_338_io_data_1_in_bits = PENetwork_37_io_to_pes_8_in_bits; // @[pe.scala 264:34]
  assign PE_338_io_data_0_in_valid = PENetwork_8_io_to_pes_15_in_valid; // @[pe.scala 264:34]
  assign PE_338_io_data_0_in_bits = PENetwork_8_io_to_pes_15_in_bits; // @[pe.scala 264:34]
  assign PE_339_clock = clock;
  assign PE_339_reset = reset;
  assign PE_339_io_data_2_sig_stat2trans = PENetwork_67_io_to_pes_9_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_339_io_data_1_in_valid = PENetwork_37_io_to_pes_9_in_valid; // @[pe.scala 264:34]
  assign PE_339_io_data_1_in_bits = PENetwork_37_io_to_pes_9_in_bits; // @[pe.scala 264:34]
  assign PE_339_io_data_0_in_valid = PENetwork_9_io_to_pes_15_in_valid; // @[pe.scala 264:34]
  assign PE_339_io_data_0_in_bits = PENetwork_9_io_to_pes_15_in_bits; // @[pe.scala 264:34]
  assign PE_340_clock = clock;
  assign PE_340_reset = reset;
  assign PE_340_io_data_2_sig_stat2trans = PENetwork_67_io_to_pes_10_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_340_io_data_1_in_valid = PENetwork_37_io_to_pes_10_in_valid; // @[pe.scala 264:34]
  assign PE_340_io_data_1_in_bits = PENetwork_37_io_to_pes_10_in_bits; // @[pe.scala 264:34]
  assign PE_340_io_data_0_in_valid = PENetwork_10_io_to_pes_15_in_valid; // @[pe.scala 264:34]
  assign PE_340_io_data_0_in_bits = PENetwork_10_io_to_pes_15_in_bits; // @[pe.scala 264:34]
  assign PE_341_clock = clock;
  assign PE_341_reset = reset;
  assign PE_341_io_data_2_sig_stat2trans = PENetwork_67_io_to_pes_11_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_341_io_data_1_in_valid = PENetwork_37_io_to_pes_11_in_valid; // @[pe.scala 264:34]
  assign PE_341_io_data_1_in_bits = PENetwork_37_io_to_pes_11_in_bits; // @[pe.scala 264:34]
  assign PE_341_io_data_0_in_valid = PENetwork_11_io_to_pes_15_in_valid; // @[pe.scala 264:34]
  assign PE_341_io_data_0_in_bits = PENetwork_11_io_to_pes_15_in_bits; // @[pe.scala 264:34]
  assign PE_342_clock = clock;
  assign PE_342_reset = reset;
  assign PE_342_io_data_2_sig_stat2trans = PENetwork_67_io_to_pes_12_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_342_io_data_1_in_valid = PENetwork_37_io_to_pes_12_in_valid; // @[pe.scala 264:34]
  assign PE_342_io_data_1_in_bits = PENetwork_37_io_to_pes_12_in_bits; // @[pe.scala 264:34]
  assign PE_342_io_data_0_in_valid = PENetwork_12_io_to_pes_15_in_valid; // @[pe.scala 264:34]
  assign PE_342_io_data_0_in_bits = PENetwork_12_io_to_pes_15_in_bits; // @[pe.scala 264:34]
  assign PE_343_clock = clock;
  assign PE_343_reset = reset;
  assign PE_343_io_data_2_sig_stat2trans = PENetwork_67_io_to_pes_13_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_343_io_data_1_in_valid = PENetwork_37_io_to_pes_13_in_valid; // @[pe.scala 264:34]
  assign PE_343_io_data_1_in_bits = PENetwork_37_io_to_pes_13_in_bits; // @[pe.scala 264:34]
  assign PE_343_io_data_0_in_valid = PENetwork_13_io_to_pes_15_in_valid; // @[pe.scala 264:34]
  assign PE_343_io_data_0_in_bits = PENetwork_13_io_to_pes_15_in_bits; // @[pe.scala 264:34]
  assign PE_344_clock = clock;
  assign PE_344_reset = reset;
  assign PE_344_io_data_2_sig_stat2trans = PENetwork_67_io_to_pes_14_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_344_io_data_1_in_valid = PENetwork_37_io_to_pes_14_in_valid; // @[pe.scala 264:34]
  assign PE_344_io_data_1_in_bits = PENetwork_37_io_to_pes_14_in_bits; // @[pe.scala 264:34]
  assign PE_344_io_data_0_in_valid = PENetwork_14_io_to_pes_15_in_valid; // @[pe.scala 264:34]
  assign PE_344_io_data_0_in_bits = PENetwork_14_io_to_pes_15_in_bits; // @[pe.scala 264:34]
  assign PE_345_clock = clock;
  assign PE_345_reset = reset;
  assign PE_345_io_data_2_sig_stat2trans = PENetwork_67_io_to_pes_15_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_345_io_data_1_in_valid = PENetwork_37_io_to_pes_15_in_valid; // @[pe.scala 264:34]
  assign PE_345_io_data_1_in_bits = PENetwork_37_io_to_pes_15_in_bits; // @[pe.scala 264:34]
  assign PE_345_io_data_0_in_valid = PENetwork_15_io_to_pes_15_in_valid; // @[pe.scala 264:34]
  assign PE_345_io_data_0_in_bits = PENetwork_15_io_to_pes_15_in_bits; // @[pe.scala 264:34]
  assign PE_346_clock = clock;
  assign PE_346_reset = reset;
  assign PE_346_io_data_2_sig_stat2trans = PENetwork_67_io_to_pes_16_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_346_io_data_1_in_valid = PENetwork_37_io_to_pes_16_in_valid; // @[pe.scala 264:34]
  assign PE_346_io_data_1_in_bits = PENetwork_37_io_to_pes_16_in_bits; // @[pe.scala 264:34]
  assign PE_346_io_data_0_in_valid = PENetwork_16_io_to_pes_15_in_valid; // @[pe.scala 264:34]
  assign PE_346_io_data_0_in_bits = PENetwork_16_io_to_pes_15_in_bits; // @[pe.scala 264:34]
  assign PE_347_clock = clock;
  assign PE_347_reset = reset;
  assign PE_347_io_data_2_sig_stat2trans = PENetwork_67_io_to_pes_17_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_347_io_data_1_in_valid = PENetwork_37_io_to_pes_17_in_valid; // @[pe.scala 264:34]
  assign PE_347_io_data_1_in_bits = PENetwork_37_io_to_pes_17_in_bits; // @[pe.scala 264:34]
  assign PE_347_io_data_0_in_valid = PENetwork_17_io_to_pes_15_in_valid; // @[pe.scala 264:34]
  assign PE_347_io_data_0_in_bits = PENetwork_17_io_to_pes_15_in_bits; // @[pe.scala 264:34]
  assign PE_348_clock = clock;
  assign PE_348_reset = reset;
  assign PE_348_io_data_2_sig_stat2trans = PENetwork_67_io_to_pes_18_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_348_io_data_1_in_valid = PENetwork_37_io_to_pes_18_in_valid; // @[pe.scala 264:34]
  assign PE_348_io_data_1_in_bits = PENetwork_37_io_to_pes_18_in_bits; // @[pe.scala 264:34]
  assign PE_348_io_data_0_in_valid = PENetwork_18_io_to_pes_15_in_valid; // @[pe.scala 264:34]
  assign PE_348_io_data_0_in_bits = PENetwork_18_io_to_pes_15_in_bits; // @[pe.scala 264:34]
  assign PE_349_clock = clock;
  assign PE_349_reset = reset;
  assign PE_349_io_data_2_sig_stat2trans = PENetwork_67_io_to_pes_19_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_349_io_data_1_in_valid = PENetwork_37_io_to_pes_19_in_valid; // @[pe.scala 264:34]
  assign PE_349_io_data_1_in_bits = PENetwork_37_io_to_pes_19_in_bits; // @[pe.scala 264:34]
  assign PE_349_io_data_0_in_valid = PENetwork_19_io_to_pes_15_in_valid; // @[pe.scala 264:34]
  assign PE_349_io_data_0_in_bits = PENetwork_19_io_to_pes_15_in_bits; // @[pe.scala 264:34]
  assign PE_350_clock = clock;
  assign PE_350_reset = reset;
  assign PE_350_io_data_2_sig_stat2trans = PENetwork_67_io_to_pes_20_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_350_io_data_1_in_valid = PENetwork_37_io_to_pes_20_in_valid; // @[pe.scala 264:34]
  assign PE_350_io_data_1_in_bits = PENetwork_37_io_to_pes_20_in_bits; // @[pe.scala 264:34]
  assign PE_350_io_data_0_in_valid = PENetwork_20_io_to_pes_15_in_valid; // @[pe.scala 264:34]
  assign PE_350_io_data_0_in_bits = PENetwork_20_io_to_pes_15_in_bits; // @[pe.scala 264:34]
  assign PE_351_clock = clock;
  assign PE_351_reset = reset;
  assign PE_351_io_data_2_sig_stat2trans = PENetwork_67_io_to_pes_21_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_351_io_data_1_in_valid = PENetwork_37_io_to_pes_21_in_valid; // @[pe.scala 264:34]
  assign PE_351_io_data_1_in_bits = PENetwork_37_io_to_pes_21_in_bits; // @[pe.scala 264:34]
  assign PE_351_io_data_0_in_valid = PENetwork_21_io_to_pes_15_in_valid; // @[pe.scala 264:34]
  assign PE_351_io_data_0_in_bits = PENetwork_21_io_to_pes_15_in_bits; // @[pe.scala 264:34]
  assign PE_352_clock = clock;
  assign PE_352_reset = reset;
  assign PE_352_io_data_2_sig_stat2trans = PENetwork_68_io_to_pes_0_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_352_io_data_1_in_valid = PENetwork_38_io_to_pes_0_in_valid; // @[pe.scala 264:34]
  assign PE_352_io_data_1_in_bits = PENetwork_38_io_to_pes_0_in_bits; // @[pe.scala 264:34]
  assign PE_352_io_data_0_in_valid = PENetwork_io_to_pes_16_in_valid; // @[pe.scala 264:34]
  assign PE_352_io_data_0_in_bits = PENetwork_io_to_pes_16_in_bits; // @[pe.scala 264:34]
  assign PE_353_clock = clock;
  assign PE_353_reset = reset;
  assign PE_353_io_data_2_sig_stat2trans = PENetwork_68_io_to_pes_1_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_353_io_data_1_in_valid = PENetwork_38_io_to_pes_1_in_valid; // @[pe.scala 264:34]
  assign PE_353_io_data_1_in_bits = PENetwork_38_io_to_pes_1_in_bits; // @[pe.scala 264:34]
  assign PE_353_io_data_0_in_valid = PENetwork_1_io_to_pes_16_in_valid; // @[pe.scala 264:34]
  assign PE_353_io_data_0_in_bits = PENetwork_1_io_to_pes_16_in_bits; // @[pe.scala 264:34]
  assign PE_354_clock = clock;
  assign PE_354_reset = reset;
  assign PE_354_io_data_2_sig_stat2trans = PENetwork_68_io_to_pes_2_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_354_io_data_1_in_valid = PENetwork_38_io_to_pes_2_in_valid; // @[pe.scala 264:34]
  assign PE_354_io_data_1_in_bits = PENetwork_38_io_to_pes_2_in_bits; // @[pe.scala 264:34]
  assign PE_354_io_data_0_in_valid = PENetwork_2_io_to_pes_16_in_valid; // @[pe.scala 264:34]
  assign PE_354_io_data_0_in_bits = PENetwork_2_io_to_pes_16_in_bits; // @[pe.scala 264:34]
  assign PE_355_clock = clock;
  assign PE_355_reset = reset;
  assign PE_355_io_data_2_sig_stat2trans = PENetwork_68_io_to_pes_3_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_355_io_data_1_in_valid = PENetwork_38_io_to_pes_3_in_valid; // @[pe.scala 264:34]
  assign PE_355_io_data_1_in_bits = PENetwork_38_io_to_pes_3_in_bits; // @[pe.scala 264:34]
  assign PE_355_io_data_0_in_valid = PENetwork_3_io_to_pes_16_in_valid; // @[pe.scala 264:34]
  assign PE_355_io_data_0_in_bits = PENetwork_3_io_to_pes_16_in_bits; // @[pe.scala 264:34]
  assign PE_356_clock = clock;
  assign PE_356_reset = reset;
  assign PE_356_io_data_2_sig_stat2trans = PENetwork_68_io_to_pes_4_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_356_io_data_1_in_valid = PENetwork_38_io_to_pes_4_in_valid; // @[pe.scala 264:34]
  assign PE_356_io_data_1_in_bits = PENetwork_38_io_to_pes_4_in_bits; // @[pe.scala 264:34]
  assign PE_356_io_data_0_in_valid = PENetwork_4_io_to_pes_16_in_valid; // @[pe.scala 264:34]
  assign PE_356_io_data_0_in_bits = PENetwork_4_io_to_pes_16_in_bits; // @[pe.scala 264:34]
  assign PE_357_clock = clock;
  assign PE_357_reset = reset;
  assign PE_357_io_data_2_sig_stat2trans = PENetwork_68_io_to_pes_5_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_357_io_data_1_in_valid = PENetwork_38_io_to_pes_5_in_valid; // @[pe.scala 264:34]
  assign PE_357_io_data_1_in_bits = PENetwork_38_io_to_pes_5_in_bits; // @[pe.scala 264:34]
  assign PE_357_io_data_0_in_valid = PENetwork_5_io_to_pes_16_in_valid; // @[pe.scala 264:34]
  assign PE_357_io_data_0_in_bits = PENetwork_5_io_to_pes_16_in_bits; // @[pe.scala 264:34]
  assign PE_358_clock = clock;
  assign PE_358_reset = reset;
  assign PE_358_io_data_2_sig_stat2trans = PENetwork_68_io_to_pes_6_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_358_io_data_1_in_valid = PENetwork_38_io_to_pes_6_in_valid; // @[pe.scala 264:34]
  assign PE_358_io_data_1_in_bits = PENetwork_38_io_to_pes_6_in_bits; // @[pe.scala 264:34]
  assign PE_358_io_data_0_in_valid = PENetwork_6_io_to_pes_16_in_valid; // @[pe.scala 264:34]
  assign PE_358_io_data_0_in_bits = PENetwork_6_io_to_pes_16_in_bits; // @[pe.scala 264:34]
  assign PE_359_clock = clock;
  assign PE_359_reset = reset;
  assign PE_359_io_data_2_sig_stat2trans = PENetwork_68_io_to_pes_7_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_359_io_data_1_in_valid = PENetwork_38_io_to_pes_7_in_valid; // @[pe.scala 264:34]
  assign PE_359_io_data_1_in_bits = PENetwork_38_io_to_pes_7_in_bits; // @[pe.scala 264:34]
  assign PE_359_io_data_0_in_valid = PENetwork_7_io_to_pes_16_in_valid; // @[pe.scala 264:34]
  assign PE_359_io_data_0_in_bits = PENetwork_7_io_to_pes_16_in_bits; // @[pe.scala 264:34]
  assign PE_360_clock = clock;
  assign PE_360_reset = reset;
  assign PE_360_io_data_2_sig_stat2trans = PENetwork_68_io_to_pes_8_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_360_io_data_1_in_valid = PENetwork_38_io_to_pes_8_in_valid; // @[pe.scala 264:34]
  assign PE_360_io_data_1_in_bits = PENetwork_38_io_to_pes_8_in_bits; // @[pe.scala 264:34]
  assign PE_360_io_data_0_in_valid = PENetwork_8_io_to_pes_16_in_valid; // @[pe.scala 264:34]
  assign PE_360_io_data_0_in_bits = PENetwork_8_io_to_pes_16_in_bits; // @[pe.scala 264:34]
  assign PE_361_clock = clock;
  assign PE_361_reset = reset;
  assign PE_361_io_data_2_sig_stat2trans = PENetwork_68_io_to_pes_9_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_361_io_data_1_in_valid = PENetwork_38_io_to_pes_9_in_valid; // @[pe.scala 264:34]
  assign PE_361_io_data_1_in_bits = PENetwork_38_io_to_pes_9_in_bits; // @[pe.scala 264:34]
  assign PE_361_io_data_0_in_valid = PENetwork_9_io_to_pes_16_in_valid; // @[pe.scala 264:34]
  assign PE_361_io_data_0_in_bits = PENetwork_9_io_to_pes_16_in_bits; // @[pe.scala 264:34]
  assign PE_362_clock = clock;
  assign PE_362_reset = reset;
  assign PE_362_io_data_2_sig_stat2trans = PENetwork_68_io_to_pes_10_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_362_io_data_1_in_valid = PENetwork_38_io_to_pes_10_in_valid; // @[pe.scala 264:34]
  assign PE_362_io_data_1_in_bits = PENetwork_38_io_to_pes_10_in_bits; // @[pe.scala 264:34]
  assign PE_362_io_data_0_in_valid = PENetwork_10_io_to_pes_16_in_valid; // @[pe.scala 264:34]
  assign PE_362_io_data_0_in_bits = PENetwork_10_io_to_pes_16_in_bits; // @[pe.scala 264:34]
  assign PE_363_clock = clock;
  assign PE_363_reset = reset;
  assign PE_363_io_data_2_sig_stat2trans = PENetwork_68_io_to_pes_11_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_363_io_data_1_in_valid = PENetwork_38_io_to_pes_11_in_valid; // @[pe.scala 264:34]
  assign PE_363_io_data_1_in_bits = PENetwork_38_io_to_pes_11_in_bits; // @[pe.scala 264:34]
  assign PE_363_io_data_0_in_valid = PENetwork_11_io_to_pes_16_in_valid; // @[pe.scala 264:34]
  assign PE_363_io_data_0_in_bits = PENetwork_11_io_to_pes_16_in_bits; // @[pe.scala 264:34]
  assign PE_364_clock = clock;
  assign PE_364_reset = reset;
  assign PE_364_io_data_2_sig_stat2trans = PENetwork_68_io_to_pes_12_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_364_io_data_1_in_valid = PENetwork_38_io_to_pes_12_in_valid; // @[pe.scala 264:34]
  assign PE_364_io_data_1_in_bits = PENetwork_38_io_to_pes_12_in_bits; // @[pe.scala 264:34]
  assign PE_364_io_data_0_in_valid = PENetwork_12_io_to_pes_16_in_valid; // @[pe.scala 264:34]
  assign PE_364_io_data_0_in_bits = PENetwork_12_io_to_pes_16_in_bits; // @[pe.scala 264:34]
  assign PE_365_clock = clock;
  assign PE_365_reset = reset;
  assign PE_365_io_data_2_sig_stat2trans = PENetwork_68_io_to_pes_13_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_365_io_data_1_in_valid = PENetwork_38_io_to_pes_13_in_valid; // @[pe.scala 264:34]
  assign PE_365_io_data_1_in_bits = PENetwork_38_io_to_pes_13_in_bits; // @[pe.scala 264:34]
  assign PE_365_io_data_0_in_valid = PENetwork_13_io_to_pes_16_in_valid; // @[pe.scala 264:34]
  assign PE_365_io_data_0_in_bits = PENetwork_13_io_to_pes_16_in_bits; // @[pe.scala 264:34]
  assign PE_366_clock = clock;
  assign PE_366_reset = reset;
  assign PE_366_io_data_2_sig_stat2trans = PENetwork_68_io_to_pes_14_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_366_io_data_1_in_valid = PENetwork_38_io_to_pes_14_in_valid; // @[pe.scala 264:34]
  assign PE_366_io_data_1_in_bits = PENetwork_38_io_to_pes_14_in_bits; // @[pe.scala 264:34]
  assign PE_366_io_data_0_in_valid = PENetwork_14_io_to_pes_16_in_valid; // @[pe.scala 264:34]
  assign PE_366_io_data_0_in_bits = PENetwork_14_io_to_pes_16_in_bits; // @[pe.scala 264:34]
  assign PE_367_clock = clock;
  assign PE_367_reset = reset;
  assign PE_367_io_data_2_sig_stat2trans = PENetwork_68_io_to_pes_15_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_367_io_data_1_in_valid = PENetwork_38_io_to_pes_15_in_valid; // @[pe.scala 264:34]
  assign PE_367_io_data_1_in_bits = PENetwork_38_io_to_pes_15_in_bits; // @[pe.scala 264:34]
  assign PE_367_io_data_0_in_valid = PENetwork_15_io_to_pes_16_in_valid; // @[pe.scala 264:34]
  assign PE_367_io_data_0_in_bits = PENetwork_15_io_to_pes_16_in_bits; // @[pe.scala 264:34]
  assign PE_368_clock = clock;
  assign PE_368_reset = reset;
  assign PE_368_io_data_2_sig_stat2trans = PENetwork_68_io_to_pes_16_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_368_io_data_1_in_valid = PENetwork_38_io_to_pes_16_in_valid; // @[pe.scala 264:34]
  assign PE_368_io_data_1_in_bits = PENetwork_38_io_to_pes_16_in_bits; // @[pe.scala 264:34]
  assign PE_368_io_data_0_in_valid = PENetwork_16_io_to_pes_16_in_valid; // @[pe.scala 264:34]
  assign PE_368_io_data_0_in_bits = PENetwork_16_io_to_pes_16_in_bits; // @[pe.scala 264:34]
  assign PE_369_clock = clock;
  assign PE_369_reset = reset;
  assign PE_369_io_data_2_sig_stat2trans = PENetwork_68_io_to_pes_17_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_369_io_data_1_in_valid = PENetwork_38_io_to_pes_17_in_valid; // @[pe.scala 264:34]
  assign PE_369_io_data_1_in_bits = PENetwork_38_io_to_pes_17_in_bits; // @[pe.scala 264:34]
  assign PE_369_io_data_0_in_valid = PENetwork_17_io_to_pes_16_in_valid; // @[pe.scala 264:34]
  assign PE_369_io_data_0_in_bits = PENetwork_17_io_to_pes_16_in_bits; // @[pe.scala 264:34]
  assign PE_370_clock = clock;
  assign PE_370_reset = reset;
  assign PE_370_io_data_2_sig_stat2trans = PENetwork_68_io_to_pes_18_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_370_io_data_1_in_valid = PENetwork_38_io_to_pes_18_in_valid; // @[pe.scala 264:34]
  assign PE_370_io_data_1_in_bits = PENetwork_38_io_to_pes_18_in_bits; // @[pe.scala 264:34]
  assign PE_370_io_data_0_in_valid = PENetwork_18_io_to_pes_16_in_valid; // @[pe.scala 264:34]
  assign PE_370_io_data_0_in_bits = PENetwork_18_io_to_pes_16_in_bits; // @[pe.scala 264:34]
  assign PE_371_clock = clock;
  assign PE_371_reset = reset;
  assign PE_371_io_data_2_sig_stat2trans = PENetwork_68_io_to_pes_19_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_371_io_data_1_in_valid = PENetwork_38_io_to_pes_19_in_valid; // @[pe.scala 264:34]
  assign PE_371_io_data_1_in_bits = PENetwork_38_io_to_pes_19_in_bits; // @[pe.scala 264:34]
  assign PE_371_io_data_0_in_valid = PENetwork_19_io_to_pes_16_in_valid; // @[pe.scala 264:34]
  assign PE_371_io_data_0_in_bits = PENetwork_19_io_to_pes_16_in_bits; // @[pe.scala 264:34]
  assign PE_372_clock = clock;
  assign PE_372_reset = reset;
  assign PE_372_io_data_2_sig_stat2trans = PENetwork_68_io_to_pes_20_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_372_io_data_1_in_valid = PENetwork_38_io_to_pes_20_in_valid; // @[pe.scala 264:34]
  assign PE_372_io_data_1_in_bits = PENetwork_38_io_to_pes_20_in_bits; // @[pe.scala 264:34]
  assign PE_372_io_data_0_in_valid = PENetwork_20_io_to_pes_16_in_valid; // @[pe.scala 264:34]
  assign PE_372_io_data_0_in_bits = PENetwork_20_io_to_pes_16_in_bits; // @[pe.scala 264:34]
  assign PE_373_clock = clock;
  assign PE_373_reset = reset;
  assign PE_373_io_data_2_sig_stat2trans = PENetwork_68_io_to_pes_21_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_373_io_data_1_in_valid = PENetwork_38_io_to_pes_21_in_valid; // @[pe.scala 264:34]
  assign PE_373_io_data_1_in_bits = PENetwork_38_io_to_pes_21_in_bits; // @[pe.scala 264:34]
  assign PE_373_io_data_0_in_valid = PENetwork_21_io_to_pes_16_in_valid; // @[pe.scala 264:34]
  assign PE_373_io_data_0_in_bits = PENetwork_21_io_to_pes_16_in_bits; // @[pe.scala 264:34]
  assign PE_374_clock = clock;
  assign PE_374_reset = reset;
  assign PE_374_io_data_2_sig_stat2trans = PENetwork_69_io_to_pes_0_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_374_io_data_1_in_valid = PENetwork_39_io_to_pes_0_in_valid; // @[pe.scala 264:34]
  assign PE_374_io_data_1_in_bits = PENetwork_39_io_to_pes_0_in_bits; // @[pe.scala 264:34]
  assign PE_374_io_data_0_in_valid = PENetwork_io_to_pes_17_in_valid; // @[pe.scala 264:34]
  assign PE_374_io_data_0_in_bits = PENetwork_io_to_pes_17_in_bits; // @[pe.scala 264:34]
  assign PE_375_clock = clock;
  assign PE_375_reset = reset;
  assign PE_375_io_data_2_sig_stat2trans = PENetwork_69_io_to_pes_1_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_375_io_data_1_in_valid = PENetwork_39_io_to_pes_1_in_valid; // @[pe.scala 264:34]
  assign PE_375_io_data_1_in_bits = PENetwork_39_io_to_pes_1_in_bits; // @[pe.scala 264:34]
  assign PE_375_io_data_0_in_valid = PENetwork_1_io_to_pes_17_in_valid; // @[pe.scala 264:34]
  assign PE_375_io_data_0_in_bits = PENetwork_1_io_to_pes_17_in_bits; // @[pe.scala 264:34]
  assign PE_376_clock = clock;
  assign PE_376_reset = reset;
  assign PE_376_io_data_2_sig_stat2trans = PENetwork_69_io_to_pes_2_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_376_io_data_1_in_valid = PENetwork_39_io_to_pes_2_in_valid; // @[pe.scala 264:34]
  assign PE_376_io_data_1_in_bits = PENetwork_39_io_to_pes_2_in_bits; // @[pe.scala 264:34]
  assign PE_376_io_data_0_in_valid = PENetwork_2_io_to_pes_17_in_valid; // @[pe.scala 264:34]
  assign PE_376_io_data_0_in_bits = PENetwork_2_io_to_pes_17_in_bits; // @[pe.scala 264:34]
  assign PE_377_clock = clock;
  assign PE_377_reset = reset;
  assign PE_377_io_data_2_sig_stat2trans = PENetwork_69_io_to_pes_3_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_377_io_data_1_in_valid = PENetwork_39_io_to_pes_3_in_valid; // @[pe.scala 264:34]
  assign PE_377_io_data_1_in_bits = PENetwork_39_io_to_pes_3_in_bits; // @[pe.scala 264:34]
  assign PE_377_io_data_0_in_valid = PENetwork_3_io_to_pes_17_in_valid; // @[pe.scala 264:34]
  assign PE_377_io_data_0_in_bits = PENetwork_3_io_to_pes_17_in_bits; // @[pe.scala 264:34]
  assign PE_378_clock = clock;
  assign PE_378_reset = reset;
  assign PE_378_io_data_2_sig_stat2trans = PENetwork_69_io_to_pes_4_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_378_io_data_1_in_valid = PENetwork_39_io_to_pes_4_in_valid; // @[pe.scala 264:34]
  assign PE_378_io_data_1_in_bits = PENetwork_39_io_to_pes_4_in_bits; // @[pe.scala 264:34]
  assign PE_378_io_data_0_in_valid = PENetwork_4_io_to_pes_17_in_valid; // @[pe.scala 264:34]
  assign PE_378_io_data_0_in_bits = PENetwork_4_io_to_pes_17_in_bits; // @[pe.scala 264:34]
  assign PE_379_clock = clock;
  assign PE_379_reset = reset;
  assign PE_379_io_data_2_sig_stat2trans = PENetwork_69_io_to_pes_5_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_379_io_data_1_in_valid = PENetwork_39_io_to_pes_5_in_valid; // @[pe.scala 264:34]
  assign PE_379_io_data_1_in_bits = PENetwork_39_io_to_pes_5_in_bits; // @[pe.scala 264:34]
  assign PE_379_io_data_0_in_valid = PENetwork_5_io_to_pes_17_in_valid; // @[pe.scala 264:34]
  assign PE_379_io_data_0_in_bits = PENetwork_5_io_to_pes_17_in_bits; // @[pe.scala 264:34]
  assign PE_380_clock = clock;
  assign PE_380_reset = reset;
  assign PE_380_io_data_2_sig_stat2trans = PENetwork_69_io_to_pes_6_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_380_io_data_1_in_valid = PENetwork_39_io_to_pes_6_in_valid; // @[pe.scala 264:34]
  assign PE_380_io_data_1_in_bits = PENetwork_39_io_to_pes_6_in_bits; // @[pe.scala 264:34]
  assign PE_380_io_data_0_in_valid = PENetwork_6_io_to_pes_17_in_valid; // @[pe.scala 264:34]
  assign PE_380_io_data_0_in_bits = PENetwork_6_io_to_pes_17_in_bits; // @[pe.scala 264:34]
  assign PE_381_clock = clock;
  assign PE_381_reset = reset;
  assign PE_381_io_data_2_sig_stat2trans = PENetwork_69_io_to_pes_7_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_381_io_data_1_in_valid = PENetwork_39_io_to_pes_7_in_valid; // @[pe.scala 264:34]
  assign PE_381_io_data_1_in_bits = PENetwork_39_io_to_pes_7_in_bits; // @[pe.scala 264:34]
  assign PE_381_io_data_0_in_valid = PENetwork_7_io_to_pes_17_in_valid; // @[pe.scala 264:34]
  assign PE_381_io_data_0_in_bits = PENetwork_7_io_to_pes_17_in_bits; // @[pe.scala 264:34]
  assign PE_382_clock = clock;
  assign PE_382_reset = reset;
  assign PE_382_io_data_2_sig_stat2trans = PENetwork_69_io_to_pes_8_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_382_io_data_1_in_valid = PENetwork_39_io_to_pes_8_in_valid; // @[pe.scala 264:34]
  assign PE_382_io_data_1_in_bits = PENetwork_39_io_to_pes_8_in_bits; // @[pe.scala 264:34]
  assign PE_382_io_data_0_in_valid = PENetwork_8_io_to_pes_17_in_valid; // @[pe.scala 264:34]
  assign PE_382_io_data_0_in_bits = PENetwork_8_io_to_pes_17_in_bits; // @[pe.scala 264:34]
  assign PE_383_clock = clock;
  assign PE_383_reset = reset;
  assign PE_383_io_data_2_sig_stat2trans = PENetwork_69_io_to_pes_9_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_383_io_data_1_in_valid = PENetwork_39_io_to_pes_9_in_valid; // @[pe.scala 264:34]
  assign PE_383_io_data_1_in_bits = PENetwork_39_io_to_pes_9_in_bits; // @[pe.scala 264:34]
  assign PE_383_io_data_0_in_valid = PENetwork_9_io_to_pes_17_in_valid; // @[pe.scala 264:34]
  assign PE_383_io_data_0_in_bits = PENetwork_9_io_to_pes_17_in_bits; // @[pe.scala 264:34]
  assign PE_384_clock = clock;
  assign PE_384_reset = reset;
  assign PE_384_io_data_2_sig_stat2trans = PENetwork_69_io_to_pes_10_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_384_io_data_1_in_valid = PENetwork_39_io_to_pes_10_in_valid; // @[pe.scala 264:34]
  assign PE_384_io_data_1_in_bits = PENetwork_39_io_to_pes_10_in_bits; // @[pe.scala 264:34]
  assign PE_384_io_data_0_in_valid = PENetwork_10_io_to_pes_17_in_valid; // @[pe.scala 264:34]
  assign PE_384_io_data_0_in_bits = PENetwork_10_io_to_pes_17_in_bits; // @[pe.scala 264:34]
  assign PE_385_clock = clock;
  assign PE_385_reset = reset;
  assign PE_385_io_data_2_sig_stat2trans = PENetwork_69_io_to_pes_11_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_385_io_data_1_in_valid = PENetwork_39_io_to_pes_11_in_valid; // @[pe.scala 264:34]
  assign PE_385_io_data_1_in_bits = PENetwork_39_io_to_pes_11_in_bits; // @[pe.scala 264:34]
  assign PE_385_io_data_0_in_valid = PENetwork_11_io_to_pes_17_in_valid; // @[pe.scala 264:34]
  assign PE_385_io_data_0_in_bits = PENetwork_11_io_to_pes_17_in_bits; // @[pe.scala 264:34]
  assign PE_386_clock = clock;
  assign PE_386_reset = reset;
  assign PE_386_io_data_2_sig_stat2trans = PENetwork_69_io_to_pes_12_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_386_io_data_1_in_valid = PENetwork_39_io_to_pes_12_in_valid; // @[pe.scala 264:34]
  assign PE_386_io_data_1_in_bits = PENetwork_39_io_to_pes_12_in_bits; // @[pe.scala 264:34]
  assign PE_386_io_data_0_in_valid = PENetwork_12_io_to_pes_17_in_valid; // @[pe.scala 264:34]
  assign PE_386_io_data_0_in_bits = PENetwork_12_io_to_pes_17_in_bits; // @[pe.scala 264:34]
  assign PE_387_clock = clock;
  assign PE_387_reset = reset;
  assign PE_387_io_data_2_sig_stat2trans = PENetwork_69_io_to_pes_13_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_387_io_data_1_in_valid = PENetwork_39_io_to_pes_13_in_valid; // @[pe.scala 264:34]
  assign PE_387_io_data_1_in_bits = PENetwork_39_io_to_pes_13_in_bits; // @[pe.scala 264:34]
  assign PE_387_io_data_0_in_valid = PENetwork_13_io_to_pes_17_in_valid; // @[pe.scala 264:34]
  assign PE_387_io_data_0_in_bits = PENetwork_13_io_to_pes_17_in_bits; // @[pe.scala 264:34]
  assign PE_388_clock = clock;
  assign PE_388_reset = reset;
  assign PE_388_io_data_2_sig_stat2trans = PENetwork_69_io_to_pes_14_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_388_io_data_1_in_valid = PENetwork_39_io_to_pes_14_in_valid; // @[pe.scala 264:34]
  assign PE_388_io_data_1_in_bits = PENetwork_39_io_to_pes_14_in_bits; // @[pe.scala 264:34]
  assign PE_388_io_data_0_in_valid = PENetwork_14_io_to_pes_17_in_valid; // @[pe.scala 264:34]
  assign PE_388_io_data_0_in_bits = PENetwork_14_io_to_pes_17_in_bits; // @[pe.scala 264:34]
  assign PE_389_clock = clock;
  assign PE_389_reset = reset;
  assign PE_389_io_data_2_sig_stat2trans = PENetwork_69_io_to_pes_15_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_389_io_data_1_in_valid = PENetwork_39_io_to_pes_15_in_valid; // @[pe.scala 264:34]
  assign PE_389_io_data_1_in_bits = PENetwork_39_io_to_pes_15_in_bits; // @[pe.scala 264:34]
  assign PE_389_io_data_0_in_valid = PENetwork_15_io_to_pes_17_in_valid; // @[pe.scala 264:34]
  assign PE_389_io_data_0_in_bits = PENetwork_15_io_to_pes_17_in_bits; // @[pe.scala 264:34]
  assign PE_390_clock = clock;
  assign PE_390_reset = reset;
  assign PE_390_io_data_2_sig_stat2trans = PENetwork_69_io_to_pes_16_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_390_io_data_1_in_valid = PENetwork_39_io_to_pes_16_in_valid; // @[pe.scala 264:34]
  assign PE_390_io_data_1_in_bits = PENetwork_39_io_to_pes_16_in_bits; // @[pe.scala 264:34]
  assign PE_390_io_data_0_in_valid = PENetwork_16_io_to_pes_17_in_valid; // @[pe.scala 264:34]
  assign PE_390_io_data_0_in_bits = PENetwork_16_io_to_pes_17_in_bits; // @[pe.scala 264:34]
  assign PE_391_clock = clock;
  assign PE_391_reset = reset;
  assign PE_391_io_data_2_sig_stat2trans = PENetwork_69_io_to_pes_17_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_391_io_data_1_in_valid = PENetwork_39_io_to_pes_17_in_valid; // @[pe.scala 264:34]
  assign PE_391_io_data_1_in_bits = PENetwork_39_io_to_pes_17_in_bits; // @[pe.scala 264:34]
  assign PE_391_io_data_0_in_valid = PENetwork_17_io_to_pes_17_in_valid; // @[pe.scala 264:34]
  assign PE_391_io_data_0_in_bits = PENetwork_17_io_to_pes_17_in_bits; // @[pe.scala 264:34]
  assign PE_392_clock = clock;
  assign PE_392_reset = reset;
  assign PE_392_io_data_2_sig_stat2trans = PENetwork_69_io_to_pes_18_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_392_io_data_1_in_valid = PENetwork_39_io_to_pes_18_in_valid; // @[pe.scala 264:34]
  assign PE_392_io_data_1_in_bits = PENetwork_39_io_to_pes_18_in_bits; // @[pe.scala 264:34]
  assign PE_392_io_data_0_in_valid = PENetwork_18_io_to_pes_17_in_valid; // @[pe.scala 264:34]
  assign PE_392_io_data_0_in_bits = PENetwork_18_io_to_pes_17_in_bits; // @[pe.scala 264:34]
  assign PE_393_clock = clock;
  assign PE_393_reset = reset;
  assign PE_393_io_data_2_sig_stat2trans = PENetwork_69_io_to_pes_19_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_393_io_data_1_in_valid = PENetwork_39_io_to_pes_19_in_valid; // @[pe.scala 264:34]
  assign PE_393_io_data_1_in_bits = PENetwork_39_io_to_pes_19_in_bits; // @[pe.scala 264:34]
  assign PE_393_io_data_0_in_valid = PENetwork_19_io_to_pes_17_in_valid; // @[pe.scala 264:34]
  assign PE_393_io_data_0_in_bits = PENetwork_19_io_to_pes_17_in_bits; // @[pe.scala 264:34]
  assign PE_394_clock = clock;
  assign PE_394_reset = reset;
  assign PE_394_io_data_2_sig_stat2trans = PENetwork_69_io_to_pes_20_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_394_io_data_1_in_valid = PENetwork_39_io_to_pes_20_in_valid; // @[pe.scala 264:34]
  assign PE_394_io_data_1_in_bits = PENetwork_39_io_to_pes_20_in_bits; // @[pe.scala 264:34]
  assign PE_394_io_data_0_in_valid = PENetwork_20_io_to_pes_17_in_valid; // @[pe.scala 264:34]
  assign PE_394_io_data_0_in_bits = PENetwork_20_io_to_pes_17_in_bits; // @[pe.scala 264:34]
  assign PE_395_clock = clock;
  assign PE_395_reset = reset;
  assign PE_395_io_data_2_sig_stat2trans = PENetwork_69_io_to_pes_21_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_395_io_data_1_in_valid = PENetwork_39_io_to_pes_21_in_valid; // @[pe.scala 264:34]
  assign PE_395_io_data_1_in_bits = PENetwork_39_io_to_pes_21_in_bits; // @[pe.scala 264:34]
  assign PE_395_io_data_0_in_valid = PENetwork_21_io_to_pes_17_in_valid; // @[pe.scala 264:34]
  assign PE_395_io_data_0_in_bits = PENetwork_21_io_to_pes_17_in_bits; // @[pe.scala 264:34]
  assign PE_396_clock = clock;
  assign PE_396_reset = reset;
  assign PE_396_io_data_2_sig_stat2trans = PENetwork_70_io_to_pes_0_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_396_io_data_1_in_valid = PENetwork_40_io_to_pes_0_in_valid; // @[pe.scala 264:34]
  assign PE_396_io_data_1_in_bits = PENetwork_40_io_to_pes_0_in_bits; // @[pe.scala 264:34]
  assign PE_396_io_data_0_in_valid = PENetwork_io_to_pes_18_in_valid; // @[pe.scala 264:34]
  assign PE_396_io_data_0_in_bits = PENetwork_io_to_pes_18_in_bits; // @[pe.scala 264:34]
  assign PE_397_clock = clock;
  assign PE_397_reset = reset;
  assign PE_397_io_data_2_sig_stat2trans = PENetwork_70_io_to_pes_1_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_397_io_data_1_in_valid = PENetwork_40_io_to_pes_1_in_valid; // @[pe.scala 264:34]
  assign PE_397_io_data_1_in_bits = PENetwork_40_io_to_pes_1_in_bits; // @[pe.scala 264:34]
  assign PE_397_io_data_0_in_valid = PENetwork_1_io_to_pes_18_in_valid; // @[pe.scala 264:34]
  assign PE_397_io_data_0_in_bits = PENetwork_1_io_to_pes_18_in_bits; // @[pe.scala 264:34]
  assign PE_398_clock = clock;
  assign PE_398_reset = reset;
  assign PE_398_io_data_2_sig_stat2trans = PENetwork_70_io_to_pes_2_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_398_io_data_1_in_valid = PENetwork_40_io_to_pes_2_in_valid; // @[pe.scala 264:34]
  assign PE_398_io_data_1_in_bits = PENetwork_40_io_to_pes_2_in_bits; // @[pe.scala 264:34]
  assign PE_398_io_data_0_in_valid = PENetwork_2_io_to_pes_18_in_valid; // @[pe.scala 264:34]
  assign PE_398_io_data_0_in_bits = PENetwork_2_io_to_pes_18_in_bits; // @[pe.scala 264:34]
  assign PE_399_clock = clock;
  assign PE_399_reset = reset;
  assign PE_399_io_data_2_sig_stat2trans = PENetwork_70_io_to_pes_3_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_399_io_data_1_in_valid = PENetwork_40_io_to_pes_3_in_valid; // @[pe.scala 264:34]
  assign PE_399_io_data_1_in_bits = PENetwork_40_io_to_pes_3_in_bits; // @[pe.scala 264:34]
  assign PE_399_io_data_0_in_valid = PENetwork_3_io_to_pes_18_in_valid; // @[pe.scala 264:34]
  assign PE_399_io_data_0_in_bits = PENetwork_3_io_to_pes_18_in_bits; // @[pe.scala 264:34]
  assign PE_400_clock = clock;
  assign PE_400_reset = reset;
  assign PE_400_io_data_2_sig_stat2trans = PENetwork_70_io_to_pes_4_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_400_io_data_1_in_valid = PENetwork_40_io_to_pes_4_in_valid; // @[pe.scala 264:34]
  assign PE_400_io_data_1_in_bits = PENetwork_40_io_to_pes_4_in_bits; // @[pe.scala 264:34]
  assign PE_400_io_data_0_in_valid = PENetwork_4_io_to_pes_18_in_valid; // @[pe.scala 264:34]
  assign PE_400_io_data_0_in_bits = PENetwork_4_io_to_pes_18_in_bits; // @[pe.scala 264:34]
  assign PE_401_clock = clock;
  assign PE_401_reset = reset;
  assign PE_401_io_data_2_sig_stat2trans = PENetwork_70_io_to_pes_5_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_401_io_data_1_in_valid = PENetwork_40_io_to_pes_5_in_valid; // @[pe.scala 264:34]
  assign PE_401_io_data_1_in_bits = PENetwork_40_io_to_pes_5_in_bits; // @[pe.scala 264:34]
  assign PE_401_io_data_0_in_valid = PENetwork_5_io_to_pes_18_in_valid; // @[pe.scala 264:34]
  assign PE_401_io_data_0_in_bits = PENetwork_5_io_to_pes_18_in_bits; // @[pe.scala 264:34]
  assign PE_402_clock = clock;
  assign PE_402_reset = reset;
  assign PE_402_io_data_2_sig_stat2trans = PENetwork_70_io_to_pes_6_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_402_io_data_1_in_valid = PENetwork_40_io_to_pes_6_in_valid; // @[pe.scala 264:34]
  assign PE_402_io_data_1_in_bits = PENetwork_40_io_to_pes_6_in_bits; // @[pe.scala 264:34]
  assign PE_402_io_data_0_in_valid = PENetwork_6_io_to_pes_18_in_valid; // @[pe.scala 264:34]
  assign PE_402_io_data_0_in_bits = PENetwork_6_io_to_pes_18_in_bits; // @[pe.scala 264:34]
  assign PE_403_clock = clock;
  assign PE_403_reset = reset;
  assign PE_403_io_data_2_sig_stat2trans = PENetwork_70_io_to_pes_7_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_403_io_data_1_in_valid = PENetwork_40_io_to_pes_7_in_valid; // @[pe.scala 264:34]
  assign PE_403_io_data_1_in_bits = PENetwork_40_io_to_pes_7_in_bits; // @[pe.scala 264:34]
  assign PE_403_io_data_0_in_valid = PENetwork_7_io_to_pes_18_in_valid; // @[pe.scala 264:34]
  assign PE_403_io_data_0_in_bits = PENetwork_7_io_to_pes_18_in_bits; // @[pe.scala 264:34]
  assign PE_404_clock = clock;
  assign PE_404_reset = reset;
  assign PE_404_io_data_2_sig_stat2trans = PENetwork_70_io_to_pes_8_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_404_io_data_1_in_valid = PENetwork_40_io_to_pes_8_in_valid; // @[pe.scala 264:34]
  assign PE_404_io_data_1_in_bits = PENetwork_40_io_to_pes_8_in_bits; // @[pe.scala 264:34]
  assign PE_404_io_data_0_in_valid = PENetwork_8_io_to_pes_18_in_valid; // @[pe.scala 264:34]
  assign PE_404_io_data_0_in_bits = PENetwork_8_io_to_pes_18_in_bits; // @[pe.scala 264:34]
  assign PE_405_clock = clock;
  assign PE_405_reset = reset;
  assign PE_405_io_data_2_sig_stat2trans = PENetwork_70_io_to_pes_9_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_405_io_data_1_in_valid = PENetwork_40_io_to_pes_9_in_valid; // @[pe.scala 264:34]
  assign PE_405_io_data_1_in_bits = PENetwork_40_io_to_pes_9_in_bits; // @[pe.scala 264:34]
  assign PE_405_io_data_0_in_valid = PENetwork_9_io_to_pes_18_in_valid; // @[pe.scala 264:34]
  assign PE_405_io_data_0_in_bits = PENetwork_9_io_to_pes_18_in_bits; // @[pe.scala 264:34]
  assign PE_406_clock = clock;
  assign PE_406_reset = reset;
  assign PE_406_io_data_2_sig_stat2trans = PENetwork_70_io_to_pes_10_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_406_io_data_1_in_valid = PENetwork_40_io_to_pes_10_in_valid; // @[pe.scala 264:34]
  assign PE_406_io_data_1_in_bits = PENetwork_40_io_to_pes_10_in_bits; // @[pe.scala 264:34]
  assign PE_406_io_data_0_in_valid = PENetwork_10_io_to_pes_18_in_valid; // @[pe.scala 264:34]
  assign PE_406_io_data_0_in_bits = PENetwork_10_io_to_pes_18_in_bits; // @[pe.scala 264:34]
  assign PE_407_clock = clock;
  assign PE_407_reset = reset;
  assign PE_407_io_data_2_sig_stat2trans = PENetwork_70_io_to_pes_11_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_407_io_data_1_in_valid = PENetwork_40_io_to_pes_11_in_valid; // @[pe.scala 264:34]
  assign PE_407_io_data_1_in_bits = PENetwork_40_io_to_pes_11_in_bits; // @[pe.scala 264:34]
  assign PE_407_io_data_0_in_valid = PENetwork_11_io_to_pes_18_in_valid; // @[pe.scala 264:34]
  assign PE_407_io_data_0_in_bits = PENetwork_11_io_to_pes_18_in_bits; // @[pe.scala 264:34]
  assign PE_408_clock = clock;
  assign PE_408_reset = reset;
  assign PE_408_io_data_2_sig_stat2trans = PENetwork_70_io_to_pes_12_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_408_io_data_1_in_valid = PENetwork_40_io_to_pes_12_in_valid; // @[pe.scala 264:34]
  assign PE_408_io_data_1_in_bits = PENetwork_40_io_to_pes_12_in_bits; // @[pe.scala 264:34]
  assign PE_408_io_data_0_in_valid = PENetwork_12_io_to_pes_18_in_valid; // @[pe.scala 264:34]
  assign PE_408_io_data_0_in_bits = PENetwork_12_io_to_pes_18_in_bits; // @[pe.scala 264:34]
  assign PE_409_clock = clock;
  assign PE_409_reset = reset;
  assign PE_409_io_data_2_sig_stat2trans = PENetwork_70_io_to_pes_13_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_409_io_data_1_in_valid = PENetwork_40_io_to_pes_13_in_valid; // @[pe.scala 264:34]
  assign PE_409_io_data_1_in_bits = PENetwork_40_io_to_pes_13_in_bits; // @[pe.scala 264:34]
  assign PE_409_io_data_0_in_valid = PENetwork_13_io_to_pes_18_in_valid; // @[pe.scala 264:34]
  assign PE_409_io_data_0_in_bits = PENetwork_13_io_to_pes_18_in_bits; // @[pe.scala 264:34]
  assign PE_410_clock = clock;
  assign PE_410_reset = reset;
  assign PE_410_io_data_2_sig_stat2trans = PENetwork_70_io_to_pes_14_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_410_io_data_1_in_valid = PENetwork_40_io_to_pes_14_in_valid; // @[pe.scala 264:34]
  assign PE_410_io_data_1_in_bits = PENetwork_40_io_to_pes_14_in_bits; // @[pe.scala 264:34]
  assign PE_410_io_data_0_in_valid = PENetwork_14_io_to_pes_18_in_valid; // @[pe.scala 264:34]
  assign PE_410_io_data_0_in_bits = PENetwork_14_io_to_pes_18_in_bits; // @[pe.scala 264:34]
  assign PE_411_clock = clock;
  assign PE_411_reset = reset;
  assign PE_411_io_data_2_sig_stat2trans = PENetwork_70_io_to_pes_15_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_411_io_data_1_in_valid = PENetwork_40_io_to_pes_15_in_valid; // @[pe.scala 264:34]
  assign PE_411_io_data_1_in_bits = PENetwork_40_io_to_pes_15_in_bits; // @[pe.scala 264:34]
  assign PE_411_io_data_0_in_valid = PENetwork_15_io_to_pes_18_in_valid; // @[pe.scala 264:34]
  assign PE_411_io_data_0_in_bits = PENetwork_15_io_to_pes_18_in_bits; // @[pe.scala 264:34]
  assign PE_412_clock = clock;
  assign PE_412_reset = reset;
  assign PE_412_io_data_2_sig_stat2trans = PENetwork_70_io_to_pes_16_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_412_io_data_1_in_valid = PENetwork_40_io_to_pes_16_in_valid; // @[pe.scala 264:34]
  assign PE_412_io_data_1_in_bits = PENetwork_40_io_to_pes_16_in_bits; // @[pe.scala 264:34]
  assign PE_412_io_data_0_in_valid = PENetwork_16_io_to_pes_18_in_valid; // @[pe.scala 264:34]
  assign PE_412_io_data_0_in_bits = PENetwork_16_io_to_pes_18_in_bits; // @[pe.scala 264:34]
  assign PE_413_clock = clock;
  assign PE_413_reset = reset;
  assign PE_413_io_data_2_sig_stat2trans = PENetwork_70_io_to_pes_17_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_413_io_data_1_in_valid = PENetwork_40_io_to_pes_17_in_valid; // @[pe.scala 264:34]
  assign PE_413_io_data_1_in_bits = PENetwork_40_io_to_pes_17_in_bits; // @[pe.scala 264:34]
  assign PE_413_io_data_0_in_valid = PENetwork_17_io_to_pes_18_in_valid; // @[pe.scala 264:34]
  assign PE_413_io_data_0_in_bits = PENetwork_17_io_to_pes_18_in_bits; // @[pe.scala 264:34]
  assign PE_414_clock = clock;
  assign PE_414_reset = reset;
  assign PE_414_io_data_2_sig_stat2trans = PENetwork_70_io_to_pes_18_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_414_io_data_1_in_valid = PENetwork_40_io_to_pes_18_in_valid; // @[pe.scala 264:34]
  assign PE_414_io_data_1_in_bits = PENetwork_40_io_to_pes_18_in_bits; // @[pe.scala 264:34]
  assign PE_414_io_data_0_in_valid = PENetwork_18_io_to_pes_18_in_valid; // @[pe.scala 264:34]
  assign PE_414_io_data_0_in_bits = PENetwork_18_io_to_pes_18_in_bits; // @[pe.scala 264:34]
  assign PE_415_clock = clock;
  assign PE_415_reset = reset;
  assign PE_415_io_data_2_sig_stat2trans = PENetwork_70_io_to_pes_19_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_415_io_data_1_in_valid = PENetwork_40_io_to_pes_19_in_valid; // @[pe.scala 264:34]
  assign PE_415_io_data_1_in_bits = PENetwork_40_io_to_pes_19_in_bits; // @[pe.scala 264:34]
  assign PE_415_io_data_0_in_valid = PENetwork_19_io_to_pes_18_in_valid; // @[pe.scala 264:34]
  assign PE_415_io_data_0_in_bits = PENetwork_19_io_to_pes_18_in_bits; // @[pe.scala 264:34]
  assign PE_416_clock = clock;
  assign PE_416_reset = reset;
  assign PE_416_io_data_2_sig_stat2trans = PENetwork_70_io_to_pes_20_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_416_io_data_1_in_valid = PENetwork_40_io_to_pes_20_in_valid; // @[pe.scala 264:34]
  assign PE_416_io_data_1_in_bits = PENetwork_40_io_to_pes_20_in_bits; // @[pe.scala 264:34]
  assign PE_416_io_data_0_in_valid = PENetwork_20_io_to_pes_18_in_valid; // @[pe.scala 264:34]
  assign PE_416_io_data_0_in_bits = PENetwork_20_io_to_pes_18_in_bits; // @[pe.scala 264:34]
  assign PE_417_clock = clock;
  assign PE_417_reset = reset;
  assign PE_417_io_data_2_sig_stat2trans = PENetwork_70_io_to_pes_21_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_417_io_data_1_in_valid = PENetwork_40_io_to_pes_21_in_valid; // @[pe.scala 264:34]
  assign PE_417_io_data_1_in_bits = PENetwork_40_io_to_pes_21_in_bits; // @[pe.scala 264:34]
  assign PE_417_io_data_0_in_valid = PENetwork_21_io_to_pes_18_in_valid; // @[pe.scala 264:34]
  assign PE_417_io_data_0_in_bits = PENetwork_21_io_to_pes_18_in_bits; // @[pe.scala 264:34]
  assign PE_418_clock = clock;
  assign PE_418_reset = reset;
  assign PE_418_io_data_2_sig_stat2trans = PENetwork_71_io_to_pes_0_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_418_io_data_1_in_valid = PENetwork_41_io_to_pes_0_in_valid; // @[pe.scala 264:34]
  assign PE_418_io_data_1_in_bits = PENetwork_41_io_to_pes_0_in_bits; // @[pe.scala 264:34]
  assign PE_418_io_data_0_in_valid = PENetwork_io_to_pes_19_in_valid; // @[pe.scala 264:34]
  assign PE_418_io_data_0_in_bits = PENetwork_io_to_pes_19_in_bits; // @[pe.scala 264:34]
  assign PE_419_clock = clock;
  assign PE_419_reset = reset;
  assign PE_419_io_data_2_sig_stat2trans = PENetwork_71_io_to_pes_1_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_419_io_data_1_in_valid = PENetwork_41_io_to_pes_1_in_valid; // @[pe.scala 264:34]
  assign PE_419_io_data_1_in_bits = PENetwork_41_io_to_pes_1_in_bits; // @[pe.scala 264:34]
  assign PE_419_io_data_0_in_valid = PENetwork_1_io_to_pes_19_in_valid; // @[pe.scala 264:34]
  assign PE_419_io_data_0_in_bits = PENetwork_1_io_to_pes_19_in_bits; // @[pe.scala 264:34]
  assign PE_420_clock = clock;
  assign PE_420_reset = reset;
  assign PE_420_io_data_2_sig_stat2trans = PENetwork_71_io_to_pes_2_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_420_io_data_1_in_valid = PENetwork_41_io_to_pes_2_in_valid; // @[pe.scala 264:34]
  assign PE_420_io_data_1_in_bits = PENetwork_41_io_to_pes_2_in_bits; // @[pe.scala 264:34]
  assign PE_420_io_data_0_in_valid = PENetwork_2_io_to_pes_19_in_valid; // @[pe.scala 264:34]
  assign PE_420_io_data_0_in_bits = PENetwork_2_io_to_pes_19_in_bits; // @[pe.scala 264:34]
  assign PE_421_clock = clock;
  assign PE_421_reset = reset;
  assign PE_421_io_data_2_sig_stat2trans = PENetwork_71_io_to_pes_3_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_421_io_data_1_in_valid = PENetwork_41_io_to_pes_3_in_valid; // @[pe.scala 264:34]
  assign PE_421_io_data_1_in_bits = PENetwork_41_io_to_pes_3_in_bits; // @[pe.scala 264:34]
  assign PE_421_io_data_0_in_valid = PENetwork_3_io_to_pes_19_in_valid; // @[pe.scala 264:34]
  assign PE_421_io_data_0_in_bits = PENetwork_3_io_to_pes_19_in_bits; // @[pe.scala 264:34]
  assign PE_422_clock = clock;
  assign PE_422_reset = reset;
  assign PE_422_io_data_2_sig_stat2trans = PENetwork_71_io_to_pes_4_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_422_io_data_1_in_valid = PENetwork_41_io_to_pes_4_in_valid; // @[pe.scala 264:34]
  assign PE_422_io_data_1_in_bits = PENetwork_41_io_to_pes_4_in_bits; // @[pe.scala 264:34]
  assign PE_422_io_data_0_in_valid = PENetwork_4_io_to_pes_19_in_valid; // @[pe.scala 264:34]
  assign PE_422_io_data_0_in_bits = PENetwork_4_io_to_pes_19_in_bits; // @[pe.scala 264:34]
  assign PE_423_clock = clock;
  assign PE_423_reset = reset;
  assign PE_423_io_data_2_sig_stat2trans = PENetwork_71_io_to_pes_5_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_423_io_data_1_in_valid = PENetwork_41_io_to_pes_5_in_valid; // @[pe.scala 264:34]
  assign PE_423_io_data_1_in_bits = PENetwork_41_io_to_pes_5_in_bits; // @[pe.scala 264:34]
  assign PE_423_io_data_0_in_valid = PENetwork_5_io_to_pes_19_in_valid; // @[pe.scala 264:34]
  assign PE_423_io_data_0_in_bits = PENetwork_5_io_to_pes_19_in_bits; // @[pe.scala 264:34]
  assign PE_424_clock = clock;
  assign PE_424_reset = reset;
  assign PE_424_io_data_2_sig_stat2trans = PENetwork_71_io_to_pes_6_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_424_io_data_1_in_valid = PENetwork_41_io_to_pes_6_in_valid; // @[pe.scala 264:34]
  assign PE_424_io_data_1_in_bits = PENetwork_41_io_to_pes_6_in_bits; // @[pe.scala 264:34]
  assign PE_424_io_data_0_in_valid = PENetwork_6_io_to_pes_19_in_valid; // @[pe.scala 264:34]
  assign PE_424_io_data_0_in_bits = PENetwork_6_io_to_pes_19_in_bits; // @[pe.scala 264:34]
  assign PE_425_clock = clock;
  assign PE_425_reset = reset;
  assign PE_425_io_data_2_sig_stat2trans = PENetwork_71_io_to_pes_7_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_425_io_data_1_in_valid = PENetwork_41_io_to_pes_7_in_valid; // @[pe.scala 264:34]
  assign PE_425_io_data_1_in_bits = PENetwork_41_io_to_pes_7_in_bits; // @[pe.scala 264:34]
  assign PE_425_io_data_0_in_valid = PENetwork_7_io_to_pes_19_in_valid; // @[pe.scala 264:34]
  assign PE_425_io_data_0_in_bits = PENetwork_7_io_to_pes_19_in_bits; // @[pe.scala 264:34]
  assign PE_426_clock = clock;
  assign PE_426_reset = reset;
  assign PE_426_io_data_2_sig_stat2trans = PENetwork_71_io_to_pes_8_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_426_io_data_1_in_valid = PENetwork_41_io_to_pes_8_in_valid; // @[pe.scala 264:34]
  assign PE_426_io_data_1_in_bits = PENetwork_41_io_to_pes_8_in_bits; // @[pe.scala 264:34]
  assign PE_426_io_data_0_in_valid = PENetwork_8_io_to_pes_19_in_valid; // @[pe.scala 264:34]
  assign PE_426_io_data_0_in_bits = PENetwork_8_io_to_pes_19_in_bits; // @[pe.scala 264:34]
  assign PE_427_clock = clock;
  assign PE_427_reset = reset;
  assign PE_427_io_data_2_sig_stat2trans = PENetwork_71_io_to_pes_9_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_427_io_data_1_in_valid = PENetwork_41_io_to_pes_9_in_valid; // @[pe.scala 264:34]
  assign PE_427_io_data_1_in_bits = PENetwork_41_io_to_pes_9_in_bits; // @[pe.scala 264:34]
  assign PE_427_io_data_0_in_valid = PENetwork_9_io_to_pes_19_in_valid; // @[pe.scala 264:34]
  assign PE_427_io_data_0_in_bits = PENetwork_9_io_to_pes_19_in_bits; // @[pe.scala 264:34]
  assign PE_428_clock = clock;
  assign PE_428_reset = reset;
  assign PE_428_io_data_2_sig_stat2trans = PENetwork_71_io_to_pes_10_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_428_io_data_1_in_valid = PENetwork_41_io_to_pes_10_in_valid; // @[pe.scala 264:34]
  assign PE_428_io_data_1_in_bits = PENetwork_41_io_to_pes_10_in_bits; // @[pe.scala 264:34]
  assign PE_428_io_data_0_in_valid = PENetwork_10_io_to_pes_19_in_valid; // @[pe.scala 264:34]
  assign PE_428_io_data_0_in_bits = PENetwork_10_io_to_pes_19_in_bits; // @[pe.scala 264:34]
  assign PE_429_clock = clock;
  assign PE_429_reset = reset;
  assign PE_429_io_data_2_sig_stat2trans = PENetwork_71_io_to_pes_11_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_429_io_data_1_in_valid = PENetwork_41_io_to_pes_11_in_valid; // @[pe.scala 264:34]
  assign PE_429_io_data_1_in_bits = PENetwork_41_io_to_pes_11_in_bits; // @[pe.scala 264:34]
  assign PE_429_io_data_0_in_valid = PENetwork_11_io_to_pes_19_in_valid; // @[pe.scala 264:34]
  assign PE_429_io_data_0_in_bits = PENetwork_11_io_to_pes_19_in_bits; // @[pe.scala 264:34]
  assign PE_430_clock = clock;
  assign PE_430_reset = reset;
  assign PE_430_io_data_2_sig_stat2trans = PENetwork_71_io_to_pes_12_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_430_io_data_1_in_valid = PENetwork_41_io_to_pes_12_in_valid; // @[pe.scala 264:34]
  assign PE_430_io_data_1_in_bits = PENetwork_41_io_to_pes_12_in_bits; // @[pe.scala 264:34]
  assign PE_430_io_data_0_in_valid = PENetwork_12_io_to_pes_19_in_valid; // @[pe.scala 264:34]
  assign PE_430_io_data_0_in_bits = PENetwork_12_io_to_pes_19_in_bits; // @[pe.scala 264:34]
  assign PE_431_clock = clock;
  assign PE_431_reset = reset;
  assign PE_431_io_data_2_sig_stat2trans = PENetwork_71_io_to_pes_13_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_431_io_data_1_in_valid = PENetwork_41_io_to_pes_13_in_valid; // @[pe.scala 264:34]
  assign PE_431_io_data_1_in_bits = PENetwork_41_io_to_pes_13_in_bits; // @[pe.scala 264:34]
  assign PE_431_io_data_0_in_valid = PENetwork_13_io_to_pes_19_in_valid; // @[pe.scala 264:34]
  assign PE_431_io_data_0_in_bits = PENetwork_13_io_to_pes_19_in_bits; // @[pe.scala 264:34]
  assign PE_432_clock = clock;
  assign PE_432_reset = reset;
  assign PE_432_io_data_2_sig_stat2trans = PENetwork_71_io_to_pes_14_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_432_io_data_1_in_valid = PENetwork_41_io_to_pes_14_in_valid; // @[pe.scala 264:34]
  assign PE_432_io_data_1_in_bits = PENetwork_41_io_to_pes_14_in_bits; // @[pe.scala 264:34]
  assign PE_432_io_data_0_in_valid = PENetwork_14_io_to_pes_19_in_valid; // @[pe.scala 264:34]
  assign PE_432_io_data_0_in_bits = PENetwork_14_io_to_pes_19_in_bits; // @[pe.scala 264:34]
  assign PE_433_clock = clock;
  assign PE_433_reset = reset;
  assign PE_433_io_data_2_sig_stat2trans = PENetwork_71_io_to_pes_15_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_433_io_data_1_in_valid = PENetwork_41_io_to_pes_15_in_valid; // @[pe.scala 264:34]
  assign PE_433_io_data_1_in_bits = PENetwork_41_io_to_pes_15_in_bits; // @[pe.scala 264:34]
  assign PE_433_io_data_0_in_valid = PENetwork_15_io_to_pes_19_in_valid; // @[pe.scala 264:34]
  assign PE_433_io_data_0_in_bits = PENetwork_15_io_to_pes_19_in_bits; // @[pe.scala 264:34]
  assign PE_434_clock = clock;
  assign PE_434_reset = reset;
  assign PE_434_io_data_2_sig_stat2trans = PENetwork_71_io_to_pes_16_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_434_io_data_1_in_valid = PENetwork_41_io_to_pes_16_in_valid; // @[pe.scala 264:34]
  assign PE_434_io_data_1_in_bits = PENetwork_41_io_to_pes_16_in_bits; // @[pe.scala 264:34]
  assign PE_434_io_data_0_in_valid = PENetwork_16_io_to_pes_19_in_valid; // @[pe.scala 264:34]
  assign PE_434_io_data_0_in_bits = PENetwork_16_io_to_pes_19_in_bits; // @[pe.scala 264:34]
  assign PE_435_clock = clock;
  assign PE_435_reset = reset;
  assign PE_435_io_data_2_sig_stat2trans = PENetwork_71_io_to_pes_17_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_435_io_data_1_in_valid = PENetwork_41_io_to_pes_17_in_valid; // @[pe.scala 264:34]
  assign PE_435_io_data_1_in_bits = PENetwork_41_io_to_pes_17_in_bits; // @[pe.scala 264:34]
  assign PE_435_io_data_0_in_valid = PENetwork_17_io_to_pes_19_in_valid; // @[pe.scala 264:34]
  assign PE_435_io_data_0_in_bits = PENetwork_17_io_to_pes_19_in_bits; // @[pe.scala 264:34]
  assign PE_436_clock = clock;
  assign PE_436_reset = reset;
  assign PE_436_io_data_2_sig_stat2trans = PENetwork_71_io_to_pes_18_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_436_io_data_1_in_valid = PENetwork_41_io_to_pes_18_in_valid; // @[pe.scala 264:34]
  assign PE_436_io_data_1_in_bits = PENetwork_41_io_to_pes_18_in_bits; // @[pe.scala 264:34]
  assign PE_436_io_data_0_in_valid = PENetwork_18_io_to_pes_19_in_valid; // @[pe.scala 264:34]
  assign PE_436_io_data_0_in_bits = PENetwork_18_io_to_pes_19_in_bits; // @[pe.scala 264:34]
  assign PE_437_clock = clock;
  assign PE_437_reset = reset;
  assign PE_437_io_data_2_sig_stat2trans = PENetwork_71_io_to_pes_19_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_437_io_data_1_in_valid = PENetwork_41_io_to_pes_19_in_valid; // @[pe.scala 264:34]
  assign PE_437_io_data_1_in_bits = PENetwork_41_io_to_pes_19_in_bits; // @[pe.scala 264:34]
  assign PE_437_io_data_0_in_valid = PENetwork_19_io_to_pes_19_in_valid; // @[pe.scala 264:34]
  assign PE_437_io_data_0_in_bits = PENetwork_19_io_to_pes_19_in_bits; // @[pe.scala 264:34]
  assign PE_438_clock = clock;
  assign PE_438_reset = reset;
  assign PE_438_io_data_2_sig_stat2trans = PENetwork_71_io_to_pes_20_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_438_io_data_1_in_valid = PENetwork_41_io_to_pes_20_in_valid; // @[pe.scala 264:34]
  assign PE_438_io_data_1_in_bits = PENetwork_41_io_to_pes_20_in_bits; // @[pe.scala 264:34]
  assign PE_438_io_data_0_in_valid = PENetwork_20_io_to_pes_19_in_valid; // @[pe.scala 264:34]
  assign PE_438_io_data_0_in_bits = PENetwork_20_io_to_pes_19_in_bits; // @[pe.scala 264:34]
  assign PE_439_clock = clock;
  assign PE_439_reset = reset;
  assign PE_439_io_data_2_sig_stat2trans = PENetwork_71_io_to_pes_21_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_439_io_data_1_in_valid = PENetwork_41_io_to_pes_21_in_valid; // @[pe.scala 264:34]
  assign PE_439_io_data_1_in_bits = PENetwork_41_io_to_pes_21_in_bits; // @[pe.scala 264:34]
  assign PE_439_io_data_0_in_valid = PENetwork_21_io_to_pes_19_in_valid; // @[pe.scala 264:34]
  assign PE_439_io_data_0_in_bits = PENetwork_21_io_to_pes_19_in_bits; // @[pe.scala 264:34]
  assign PE_440_clock = clock;
  assign PE_440_reset = reset;
  assign PE_440_io_data_2_sig_stat2trans = PENetwork_72_io_to_pes_0_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_440_io_data_1_in_valid = PENetwork_42_io_to_pes_0_in_valid; // @[pe.scala 264:34]
  assign PE_440_io_data_1_in_bits = PENetwork_42_io_to_pes_0_in_bits; // @[pe.scala 264:34]
  assign PE_440_io_data_0_in_valid = PENetwork_io_to_pes_20_in_valid; // @[pe.scala 264:34]
  assign PE_440_io_data_0_in_bits = PENetwork_io_to_pes_20_in_bits; // @[pe.scala 264:34]
  assign PE_441_clock = clock;
  assign PE_441_reset = reset;
  assign PE_441_io_data_2_sig_stat2trans = PENetwork_72_io_to_pes_1_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_441_io_data_1_in_valid = PENetwork_42_io_to_pes_1_in_valid; // @[pe.scala 264:34]
  assign PE_441_io_data_1_in_bits = PENetwork_42_io_to_pes_1_in_bits; // @[pe.scala 264:34]
  assign PE_441_io_data_0_in_valid = PENetwork_1_io_to_pes_20_in_valid; // @[pe.scala 264:34]
  assign PE_441_io_data_0_in_bits = PENetwork_1_io_to_pes_20_in_bits; // @[pe.scala 264:34]
  assign PE_442_clock = clock;
  assign PE_442_reset = reset;
  assign PE_442_io_data_2_sig_stat2trans = PENetwork_72_io_to_pes_2_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_442_io_data_1_in_valid = PENetwork_42_io_to_pes_2_in_valid; // @[pe.scala 264:34]
  assign PE_442_io_data_1_in_bits = PENetwork_42_io_to_pes_2_in_bits; // @[pe.scala 264:34]
  assign PE_442_io_data_0_in_valid = PENetwork_2_io_to_pes_20_in_valid; // @[pe.scala 264:34]
  assign PE_442_io_data_0_in_bits = PENetwork_2_io_to_pes_20_in_bits; // @[pe.scala 264:34]
  assign PE_443_clock = clock;
  assign PE_443_reset = reset;
  assign PE_443_io_data_2_sig_stat2trans = PENetwork_72_io_to_pes_3_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_443_io_data_1_in_valid = PENetwork_42_io_to_pes_3_in_valid; // @[pe.scala 264:34]
  assign PE_443_io_data_1_in_bits = PENetwork_42_io_to_pes_3_in_bits; // @[pe.scala 264:34]
  assign PE_443_io_data_0_in_valid = PENetwork_3_io_to_pes_20_in_valid; // @[pe.scala 264:34]
  assign PE_443_io_data_0_in_bits = PENetwork_3_io_to_pes_20_in_bits; // @[pe.scala 264:34]
  assign PE_444_clock = clock;
  assign PE_444_reset = reset;
  assign PE_444_io_data_2_sig_stat2trans = PENetwork_72_io_to_pes_4_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_444_io_data_1_in_valid = PENetwork_42_io_to_pes_4_in_valid; // @[pe.scala 264:34]
  assign PE_444_io_data_1_in_bits = PENetwork_42_io_to_pes_4_in_bits; // @[pe.scala 264:34]
  assign PE_444_io_data_0_in_valid = PENetwork_4_io_to_pes_20_in_valid; // @[pe.scala 264:34]
  assign PE_444_io_data_0_in_bits = PENetwork_4_io_to_pes_20_in_bits; // @[pe.scala 264:34]
  assign PE_445_clock = clock;
  assign PE_445_reset = reset;
  assign PE_445_io_data_2_sig_stat2trans = PENetwork_72_io_to_pes_5_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_445_io_data_1_in_valid = PENetwork_42_io_to_pes_5_in_valid; // @[pe.scala 264:34]
  assign PE_445_io_data_1_in_bits = PENetwork_42_io_to_pes_5_in_bits; // @[pe.scala 264:34]
  assign PE_445_io_data_0_in_valid = PENetwork_5_io_to_pes_20_in_valid; // @[pe.scala 264:34]
  assign PE_445_io_data_0_in_bits = PENetwork_5_io_to_pes_20_in_bits; // @[pe.scala 264:34]
  assign PE_446_clock = clock;
  assign PE_446_reset = reset;
  assign PE_446_io_data_2_sig_stat2trans = PENetwork_72_io_to_pes_6_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_446_io_data_1_in_valid = PENetwork_42_io_to_pes_6_in_valid; // @[pe.scala 264:34]
  assign PE_446_io_data_1_in_bits = PENetwork_42_io_to_pes_6_in_bits; // @[pe.scala 264:34]
  assign PE_446_io_data_0_in_valid = PENetwork_6_io_to_pes_20_in_valid; // @[pe.scala 264:34]
  assign PE_446_io_data_0_in_bits = PENetwork_6_io_to_pes_20_in_bits; // @[pe.scala 264:34]
  assign PE_447_clock = clock;
  assign PE_447_reset = reset;
  assign PE_447_io_data_2_sig_stat2trans = PENetwork_72_io_to_pes_7_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_447_io_data_1_in_valid = PENetwork_42_io_to_pes_7_in_valid; // @[pe.scala 264:34]
  assign PE_447_io_data_1_in_bits = PENetwork_42_io_to_pes_7_in_bits; // @[pe.scala 264:34]
  assign PE_447_io_data_0_in_valid = PENetwork_7_io_to_pes_20_in_valid; // @[pe.scala 264:34]
  assign PE_447_io_data_0_in_bits = PENetwork_7_io_to_pes_20_in_bits; // @[pe.scala 264:34]
  assign PE_448_clock = clock;
  assign PE_448_reset = reset;
  assign PE_448_io_data_2_sig_stat2trans = PENetwork_72_io_to_pes_8_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_448_io_data_1_in_valid = PENetwork_42_io_to_pes_8_in_valid; // @[pe.scala 264:34]
  assign PE_448_io_data_1_in_bits = PENetwork_42_io_to_pes_8_in_bits; // @[pe.scala 264:34]
  assign PE_448_io_data_0_in_valid = PENetwork_8_io_to_pes_20_in_valid; // @[pe.scala 264:34]
  assign PE_448_io_data_0_in_bits = PENetwork_8_io_to_pes_20_in_bits; // @[pe.scala 264:34]
  assign PE_449_clock = clock;
  assign PE_449_reset = reset;
  assign PE_449_io_data_2_sig_stat2trans = PENetwork_72_io_to_pes_9_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_449_io_data_1_in_valid = PENetwork_42_io_to_pes_9_in_valid; // @[pe.scala 264:34]
  assign PE_449_io_data_1_in_bits = PENetwork_42_io_to_pes_9_in_bits; // @[pe.scala 264:34]
  assign PE_449_io_data_0_in_valid = PENetwork_9_io_to_pes_20_in_valid; // @[pe.scala 264:34]
  assign PE_449_io_data_0_in_bits = PENetwork_9_io_to_pes_20_in_bits; // @[pe.scala 264:34]
  assign PE_450_clock = clock;
  assign PE_450_reset = reset;
  assign PE_450_io_data_2_sig_stat2trans = PENetwork_72_io_to_pes_10_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_450_io_data_1_in_valid = PENetwork_42_io_to_pes_10_in_valid; // @[pe.scala 264:34]
  assign PE_450_io_data_1_in_bits = PENetwork_42_io_to_pes_10_in_bits; // @[pe.scala 264:34]
  assign PE_450_io_data_0_in_valid = PENetwork_10_io_to_pes_20_in_valid; // @[pe.scala 264:34]
  assign PE_450_io_data_0_in_bits = PENetwork_10_io_to_pes_20_in_bits; // @[pe.scala 264:34]
  assign PE_451_clock = clock;
  assign PE_451_reset = reset;
  assign PE_451_io_data_2_sig_stat2trans = PENetwork_72_io_to_pes_11_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_451_io_data_1_in_valid = PENetwork_42_io_to_pes_11_in_valid; // @[pe.scala 264:34]
  assign PE_451_io_data_1_in_bits = PENetwork_42_io_to_pes_11_in_bits; // @[pe.scala 264:34]
  assign PE_451_io_data_0_in_valid = PENetwork_11_io_to_pes_20_in_valid; // @[pe.scala 264:34]
  assign PE_451_io_data_0_in_bits = PENetwork_11_io_to_pes_20_in_bits; // @[pe.scala 264:34]
  assign PE_452_clock = clock;
  assign PE_452_reset = reset;
  assign PE_452_io_data_2_sig_stat2trans = PENetwork_72_io_to_pes_12_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_452_io_data_1_in_valid = PENetwork_42_io_to_pes_12_in_valid; // @[pe.scala 264:34]
  assign PE_452_io_data_1_in_bits = PENetwork_42_io_to_pes_12_in_bits; // @[pe.scala 264:34]
  assign PE_452_io_data_0_in_valid = PENetwork_12_io_to_pes_20_in_valid; // @[pe.scala 264:34]
  assign PE_452_io_data_0_in_bits = PENetwork_12_io_to_pes_20_in_bits; // @[pe.scala 264:34]
  assign PE_453_clock = clock;
  assign PE_453_reset = reset;
  assign PE_453_io_data_2_sig_stat2trans = PENetwork_72_io_to_pes_13_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_453_io_data_1_in_valid = PENetwork_42_io_to_pes_13_in_valid; // @[pe.scala 264:34]
  assign PE_453_io_data_1_in_bits = PENetwork_42_io_to_pes_13_in_bits; // @[pe.scala 264:34]
  assign PE_453_io_data_0_in_valid = PENetwork_13_io_to_pes_20_in_valid; // @[pe.scala 264:34]
  assign PE_453_io_data_0_in_bits = PENetwork_13_io_to_pes_20_in_bits; // @[pe.scala 264:34]
  assign PE_454_clock = clock;
  assign PE_454_reset = reset;
  assign PE_454_io_data_2_sig_stat2trans = PENetwork_72_io_to_pes_14_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_454_io_data_1_in_valid = PENetwork_42_io_to_pes_14_in_valid; // @[pe.scala 264:34]
  assign PE_454_io_data_1_in_bits = PENetwork_42_io_to_pes_14_in_bits; // @[pe.scala 264:34]
  assign PE_454_io_data_0_in_valid = PENetwork_14_io_to_pes_20_in_valid; // @[pe.scala 264:34]
  assign PE_454_io_data_0_in_bits = PENetwork_14_io_to_pes_20_in_bits; // @[pe.scala 264:34]
  assign PE_455_clock = clock;
  assign PE_455_reset = reset;
  assign PE_455_io_data_2_sig_stat2trans = PENetwork_72_io_to_pes_15_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_455_io_data_1_in_valid = PENetwork_42_io_to_pes_15_in_valid; // @[pe.scala 264:34]
  assign PE_455_io_data_1_in_bits = PENetwork_42_io_to_pes_15_in_bits; // @[pe.scala 264:34]
  assign PE_455_io_data_0_in_valid = PENetwork_15_io_to_pes_20_in_valid; // @[pe.scala 264:34]
  assign PE_455_io_data_0_in_bits = PENetwork_15_io_to_pes_20_in_bits; // @[pe.scala 264:34]
  assign PE_456_clock = clock;
  assign PE_456_reset = reset;
  assign PE_456_io_data_2_sig_stat2trans = PENetwork_72_io_to_pes_16_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_456_io_data_1_in_valid = PENetwork_42_io_to_pes_16_in_valid; // @[pe.scala 264:34]
  assign PE_456_io_data_1_in_bits = PENetwork_42_io_to_pes_16_in_bits; // @[pe.scala 264:34]
  assign PE_456_io_data_0_in_valid = PENetwork_16_io_to_pes_20_in_valid; // @[pe.scala 264:34]
  assign PE_456_io_data_0_in_bits = PENetwork_16_io_to_pes_20_in_bits; // @[pe.scala 264:34]
  assign PE_457_clock = clock;
  assign PE_457_reset = reset;
  assign PE_457_io_data_2_sig_stat2trans = PENetwork_72_io_to_pes_17_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_457_io_data_1_in_valid = PENetwork_42_io_to_pes_17_in_valid; // @[pe.scala 264:34]
  assign PE_457_io_data_1_in_bits = PENetwork_42_io_to_pes_17_in_bits; // @[pe.scala 264:34]
  assign PE_457_io_data_0_in_valid = PENetwork_17_io_to_pes_20_in_valid; // @[pe.scala 264:34]
  assign PE_457_io_data_0_in_bits = PENetwork_17_io_to_pes_20_in_bits; // @[pe.scala 264:34]
  assign PE_458_clock = clock;
  assign PE_458_reset = reset;
  assign PE_458_io_data_2_sig_stat2trans = PENetwork_72_io_to_pes_18_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_458_io_data_1_in_valid = PENetwork_42_io_to_pes_18_in_valid; // @[pe.scala 264:34]
  assign PE_458_io_data_1_in_bits = PENetwork_42_io_to_pes_18_in_bits; // @[pe.scala 264:34]
  assign PE_458_io_data_0_in_valid = PENetwork_18_io_to_pes_20_in_valid; // @[pe.scala 264:34]
  assign PE_458_io_data_0_in_bits = PENetwork_18_io_to_pes_20_in_bits; // @[pe.scala 264:34]
  assign PE_459_clock = clock;
  assign PE_459_reset = reset;
  assign PE_459_io_data_2_sig_stat2trans = PENetwork_72_io_to_pes_19_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_459_io_data_1_in_valid = PENetwork_42_io_to_pes_19_in_valid; // @[pe.scala 264:34]
  assign PE_459_io_data_1_in_bits = PENetwork_42_io_to_pes_19_in_bits; // @[pe.scala 264:34]
  assign PE_459_io_data_0_in_valid = PENetwork_19_io_to_pes_20_in_valid; // @[pe.scala 264:34]
  assign PE_459_io_data_0_in_bits = PENetwork_19_io_to_pes_20_in_bits; // @[pe.scala 264:34]
  assign PE_460_clock = clock;
  assign PE_460_reset = reset;
  assign PE_460_io_data_2_sig_stat2trans = PENetwork_72_io_to_pes_20_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_460_io_data_1_in_valid = PENetwork_42_io_to_pes_20_in_valid; // @[pe.scala 264:34]
  assign PE_460_io_data_1_in_bits = PENetwork_42_io_to_pes_20_in_bits; // @[pe.scala 264:34]
  assign PE_460_io_data_0_in_valid = PENetwork_20_io_to_pes_20_in_valid; // @[pe.scala 264:34]
  assign PE_460_io_data_0_in_bits = PENetwork_20_io_to_pes_20_in_bits; // @[pe.scala 264:34]
  assign PE_461_clock = clock;
  assign PE_461_reset = reset;
  assign PE_461_io_data_2_sig_stat2trans = PENetwork_72_io_to_pes_21_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_461_io_data_1_in_valid = PENetwork_42_io_to_pes_21_in_valid; // @[pe.scala 264:34]
  assign PE_461_io_data_1_in_bits = PENetwork_42_io_to_pes_21_in_bits; // @[pe.scala 264:34]
  assign PE_461_io_data_0_in_valid = PENetwork_21_io_to_pes_20_in_valid; // @[pe.scala 264:34]
  assign PE_461_io_data_0_in_bits = PENetwork_21_io_to_pes_20_in_bits; // @[pe.scala 264:34]
  assign PE_462_clock = clock;
  assign PE_462_reset = reset;
  assign PE_462_io_data_2_sig_stat2trans = PENetwork_73_io_to_pes_0_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_462_io_data_1_in_valid = PENetwork_43_io_to_pes_0_in_valid; // @[pe.scala 264:34]
  assign PE_462_io_data_1_in_bits = PENetwork_43_io_to_pes_0_in_bits; // @[pe.scala 264:34]
  assign PE_462_io_data_0_in_valid = PENetwork_io_to_pes_21_in_valid; // @[pe.scala 264:34]
  assign PE_462_io_data_0_in_bits = PENetwork_io_to_pes_21_in_bits; // @[pe.scala 264:34]
  assign PE_463_clock = clock;
  assign PE_463_reset = reset;
  assign PE_463_io_data_2_sig_stat2trans = PENetwork_73_io_to_pes_1_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_463_io_data_1_in_valid = PENetwork_43_io_to_pes_1_in_valid; // @[pe.scala 264:34]
  assign PE_463_io_data_1_in_bits = PENetwork_43_io_to_pes_1_in_bits; // @[pe.scala 264:34]
  assign PE_463_io_data_0_in_valid = PENetwork_1_io_to_pes_21_in_valid; // @[pe.scala 264:34]
  assign PE_463_io_data_0_in_bits = PENetwork_1_io_to_pes_21_in_bits; // @[pe.scala 264:34]
  assign PE_464_clock = clock;
  assign PE_464_reset = reset;
  assign PE_464_io_data_2_sig_stat2trans = PENetwork_73_io_to_pes_2_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_464_io_data_1_in_valid = PENetwork_43_io_to_pes_2_in_valid; // @[pe.scala 264:34]
  assign PE_464_io_data_1_in_bits = PENetwork_43_io_to_pes_2_in_bits; // @[pe.scala 264:34]
  assign PE_464_io_data_0_in_valid = PENetwork_2_io_to_pes_21_in_valid; // @[pe.scala 264:34]
  assign PE_464_io_data_0_in_bits = PENetwork_2_io_to_pes_21_in_bits; // @[pe.scala 264:34]
  assign PE_465_clock = clock;
  assign PE_465_reset = reset;
  assign PE_465_io_data_2_sig_stat2trans = PENetwork_73_io_to_pes_3_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_465_io_data_1_in_valid = PENetwork_43_io_to_pes_3_in_valid; // @[pe.scala 264:34]
  assign PE_465_io_data_1_in_bits = PENetwork_43_io_to_pes_3_in_bits; // @[pe.scala 264:34]
  assign PE_465_io_data_0_in_valid = PENetwork_3_io_to_pes_21_in_valid; // @[pe.scala 264:34]
  assign PE_465_io_data_0_in_bits = PENetwork_3_io_to_pes_21_in_bits; // @[pe.scala 264:34]
  assign PE_466_clock = clock;
  assign PE_466_reset = reset;
  assign PE_466_io_data_2_sig_stat2trans = PENetwork_73_io_to_pes_4_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_466_io_data_1_in_valid = PENetwork_43_io_to_pes_4_in_valid; // @[pe.scala 264:34]
  assign PE_466_io_data_1_in_bits = PENetwork_43_io_to_pes_4_in_bits; // @[pe.scala 264:34]
  assign PE_466_io_data_0_in_valid = PENetwork_4_io_to_pes_21_in_valid; // @[pe.scala 264:34]
  assign PE_466_io_data_0_in_bits = PENetwork_4_io_to_pes_21_in_bits; // @[pe.scala 264:34]
  assign PE_467_clock = clock;
  assign PE_467_reset = reset;
  assign PE_467_io_data_2_sig_stat2trans = PENetwork_73_io_to_pes_5_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_467_io_data_1_in_valid = PENetwork_43_io_to_pes_5_in_valid; // @[pe.scala 264:34]
  assign PE_467_io_data_1_in_bits = PENetwork_43_io_to_pes_5_in_bits; // @[pe.scala 264:34]
  assign PE_467_io_data_0_in_valid = PENetwork_5_io_to_pes_21_in_valid; // @[pe.scala 264:34]
  assign PE_467_io_data_0_in_bits = PENetwork_5_io_to_pes_21_in_bits; // @[pe.scala 264:34]
  assign PE_468_clock = clock;
  assign PE_468_reset = reset;
  assign PE_468_io_data_2_sig_stat2trans = PENetwork_73_io_to_pes_6_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_468_io_data_1_in_valid = PENetwork_43_io_to_pes_6_in_valid; // @[pe.scala 264:34]
  assign PE_468_io_data_1_in_bits = PENetwork_43_io_to_pes_6_in_bits; // @[pe.scala 264:34]
  assign PE_468_io_data_0_in_valid = PENetwork_6_io_to_pes_21_in_valid; // @[pe.scala 264:34]
  assign PE_468_io_data_0_in_bits = PENetwork_6_io_to_pes_21_in_bits; // @[pe.scala 264:34]
  assign PE_469_clock = clock;
  assign PE_469_reset = reset;
  assign PE_469_io_data_2_sig_stat2trans = PENetwork_73_io_to_pes_7_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_469_io_data_1_in_valid = PENetwork_43_io_to_pes_7_in_valid; // @[pe.scala 264:34]
  assign PE_469_io_data_1_in_bits = PENetwork_43_io_to_pes_7_in_bits; // @[pe.scala 264:34]
  assign PE_469_io_data_0_in_valid = PENetwork_7_io_to_pes_21_in_valid; // @[pe.scala 264:34]
  assign PE_469_io_data_0_in_bits = PENetwork_7_io_to_pes_21_in_bits; // @[pe.scala 264:34]
  assign PE_470_clock = clock;
  assign PE_470_reset = reset;
  assign PE_470_io_data_2_sig_stat2trans = PENetwork_73_io_to_pes_8_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_470_io_data_1_in_valid = PENetwork_43_io_to_pes_8_in_valid; // @[pe.scala 264:34]
  assign PE_470_io_data_1_in_bits = PENetwork_43_io_to_pes_8_in_bits; // @[pe.scala 264:34]
  assign PE_470_io_data_0_in_valid = PENetwork_8_io_to_pes_21_in_valid; // @[pe.scala 264:34]
  assign PE_470_io_data_0_in_bits = PENetwork_8_io_to_pes_21_in_bits; // @[pe.scala 264:34]
  assign PE_471_clock = clock;
  assign PE_471_reset = reset;
  assign PE_471_io_data_2_sig_stat2trans = PENetwork_73_io_to_pes_9_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_471_io_data_1_in_valid = PENetwork_43_io_to_pes_9_in_valid; // @[pe.scala 264:34]
  assign PE_471_io_data_1_in_bits = PENetwork_43_io_to_pes_9_in_bits; // @[pe.scala 264:34]
  assign PE_471_io_data_0_in_valid = PENetwork_9_io_to_pes_21_in_valid; // @[pe.scala 264:34]
  assign PE_471_io_data_0_in_bits = PENetwork_9_io_to_pes_21_in_bits; // @[pe.scala 264:34]
  assign PE_472_clock = clock;
  assign PE_472_reset = reset;
  assign PE_472_io_data_2_sig_stat2trans = PENetwork_73_io_to_pes_10_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_472_io_data_1_in_valid = PENetwork_43_io_to_pes_10_in_valid; // @[pe.scala 264:34]
  assign PE_472_io_data_1_in_bits = PENetwork_43_io_to_pes_10_in_bits; // @[pe.scala 264:34]
  assign PE_472_io_data_0_in_valid = PENetwork_10_io_to_pes_21_in_valid; // @[pe.scala 264:34]
  assign PE_472_io_data_0_in_bits = PENetwork_10_io_to_pes_21_in_bits; // @[pe.scala 264:34]
  assign PE_473_clock = clock;
  assign PE_473_reset = reset;
  assign PE_473_io_data_2_sig_stat2trans = PENetwork_73_io_to_pes_11_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_473_io_data_1_in_valid = PENetwork_43_io_to_pes_11_in_valid; // @[pe.scala 264:34]
  assign PE_473_io_data_1_in_bits = PENetwork_43_io_to_pes_11_in_bits; // @[pe.scala 264:34]
  assign PE_473_io_data_0_in_valid = PENetwork_11_io_to_pes_21_in_valid; // @[pe.scala 264:34]
  assign PE_473_io_data_0_in_bits = PENetwork_11_io_to_pes_21_in_bits; // @[pe.scala 264:34]
  assign PE_474_clock = clock;
  assign PE_474_reset = reset;
  assign PE_474_io_data_2_sig_stat2trans = PENetwork_73_io_to_pes_12_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_474_io_data_1_in_valid = PENetwork_43_io_to_pes_12_in_valid; // @[pe.scala 264:34]
  assign PE_474_io_data_1_in_bits = PENetwork_43_io_to_pes_12_in_bits; // @[pe.scala 264:34]
  assign PE_474_io_data_0_in_valid = PENetwork_12_io_to_pes_21_in_valid; // @[pe.scala 264:34]
  assign PE_474_io_data_0_in_bits = PENetwork_12_io_to_pes_21_in_bits; // @[pe.scala 264:34]
  assign PE_475_clock = clock;
  assign PE_475_reset = reset;
  assign PE_475_io_data_2_sig_stat2trans = PENetwork_73_io_to_pes_13_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_475_io_data_1_in_valid = PENetwork_43_io_to_pes_13_in_valid; // @[pe.scala 264:34]
  assign PE_475_io_data_1_in_bits = PENetwork_43_io_to_pes_13_in_bits; // @[pe.scala 264:34]
  assign PE_475_io_data_0_in_valid = PENetwork_13_io_to_pes_21_in_valid; // @[pe.scala 264:34]
  assign PE_475_io_data_0_in_bits = PENetwork_13_io_to_pes_21_in_bits; // @[pe.scala 264:34]
  assign PE_476_clock = clock;
  assign PE_476_reset = reset;
  assign PE_476_io_data_2_sig_stat2trans = PENetwork_73_io_to_pes_14_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_476_io_data_1_in_valid = PENetwork_43_io_to_pes_14_in_valid; // @[pe.scala 264:34]
  assign PE_476_io_data_1_in_bits = PENetwork_43_io_to_pes_14_in_bits; // @[pe.scala 264:34]
  assign PE_476_io_data_0_in_valid = PENetwork_14_io_to_pes_21_in_valid; // @[pe.scala 264:34]
  assign PE_476_io_data_0_in_bits = PENetwork_14_io_to_pes_21_in_bits; // @[pe.scala 264:34]
  assign PE_477_clock = clock;
  assign PE_477_reset = reset;
  assign PE_477_io_data_2_sig_stat2trans = PENetwork_73_io_to_pes_15_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_477_io_data_1_in_valid = PENetwork_43_io_to_pes_15_in_valid; // @[pe.scala 264:34]
  assign PE_477_io_data_1_in_bits = PENetwork_43_io_to_pes_15_in_bits; // @[pe.scala 264:34]
  assign PE_477_io_data_0_in_valid = PENetwork_15_io_to_pes_21_in_valid; // @[pe.scala 264:34]
  assign PE_477_io_data_0_in_bits = PENetwork_15_io_to_pes_21_in_bits; // @[pe.scala 264:34]
  assign PE_478_clock = clock;
  assign PE_478_reset = reset;
  assign PE_478_io_data_2_sig_stat2trans = PENetwork_73_io_to_pes_16_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_478_io_data_1_in_valid = PENetwork_43_io_to_pes_16_in_valid; // @[pe.scala 264:34]
  assign PE_478_io_data_1_in_bits = PENetwork_43_io_to_pes_16_in_bits; // @[pe.scala 264:34]
  assign PE_478_io_data_0_in_valid = PENetwork_16_io_to_pes_21_in_valid; // @[pe.scala 264:34]
  assign PE_478_io_data_0_in_bits = PENetwork_16_io_to_pes_21_in_bits; // @[pe.scala 264:34]
  assign PE_479_clock = clock;
  assign PE_479_reset = reset;
  assign PE_479_io_data_2_sig_stat2trans = PENetwork_73_io_to_pes_17_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_479_io_data_1_in_valid = PENetwork_43_io_to_pes_17_in_valid; // @[pe.scala 264:34]
  assign PE_479_io_data_1_in_bits = PENetwork_43_io_to_pes_17_in_bits; // @[pe.scala 264:34]
  assign PE_479_io_data_0_in_valid = PENetwork_17_io_to_pes_21_in_valid; // @[pe.scala 264:34]
  assign PE_479_io_data_0_in_bits = PENetwork_17_io_to_pes_21_in_bits; // @[pe.scala 264:34]
  assign PE_480_clock = clock;
  assign PE_480_reset = reset;
  assign PE_480_io_data_2_sig_stat2trans = PENetwork_73_io_to_pes_18_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_480_io_data_1_in_valid = PENetwork_43_io_to_pes_18_in_valid; // @[pe.scala 264:34]
  assign PE_480_io_data_1_in_bits = PENetwork_43_io_to_pes_18_in_bits; // @[pe.scala 264:34]
  assign PE_480_io_data_0_in_valid = PENetwork_18_io_to_pes_21_in_valid; // @[pe.scala 264:34]
  assign PE_480_io_data_0_in_bits = PENetwork_18_io_to_pes_21_in_bits; // @[pe.scala 264:34]
  assign PE_481_clock = clock;
  assign PE_481_reset = reset;
  assign PE_481_io_data_2_sig_stat2trans = PENetwork_73_io_to_pes_19_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_481_io_data_1_in_valid = PENetwork_43_io_to_pes_19_in_valid; // @[pe.scala 264:34]
  assign PE_481_io_data_1_in_bits = PENetwork_43_io_to_pes_19_in_bits; // @[pe.scala 264:34]
  assign PE_481_io_data_0_in_valid = PENetwork_19_io_to_pes_21_in_valid; // @[pe.scala 264:34]
  assign PE_481_io_data_0_in_bits = PENetwork_19_io_to_pes_21_in_bits; // @[pe.scala 264:34]
  assign PE_482_clock = clock;
  assign PE_482_reset = reset;
  assign PE_482_io_data_2_sig_stat2trans = PENetwork_73_io_to_pes_20_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_482_io_data_1_in_valid = PENetwork_43_io_to_pes_20_in_valid; // @[pe.scala 264:34]
  assign PE_482_io_data_1_in_bits = PENetwork_43_io_to_pes_20_in_bits; // @[pe.scala 264:34]
  assign PE_482_io_data_0_in_valid = PENetwork_20_io_to_pes_21_in_valid; // @[pe.scala 264:34]
  assign PE_482_io_data_0_in_bits = PENetwork_20_io_to_pes_21_in_bits; // @[pe.scala 264:34]
  assign PE_483_clock = clock;
  assign PE_483_reset = reset;
  assign PE_483_io_data_2_sig_stat2trans = PENetwork_73_io_to_pes_21_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_483_io_data_1_in_valid = PENetwork_43_io_to_pes_21_in_valid; // @[pe.scala 264:34]
  assign PE_483_io_data_1_in_bits = PENetwork_43_io_to_pes_21_in_bits; // @[pe.scala 264:34]
  assign PE_483_io_data_0_in_valid = PENetwork_21_io_to_pes_21_in_valid; // @[pe.scala 264:34]
  assign PE_483_io_data_0_in_bits = PENetwork_21_io_to_pes_21_in_bits; // @[pe.scala 264:34]
  assign PE_484_clock = clock;
  assign PE_484_reset = reset;
  assign PE_484_io_data_2_sig_stat2trans = PENetwork_74_io_to_pes_0_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_484_io_data_1_in_valid = PENetwork_44_io_to_pes_0_in_valid; // @[pe.scala 264:34]
  assign PE_484_io_data_1_in_bits = PENetwork_44_io_to_pes_0_in_bits; // @[pe.scala 264:34]
  assign PE_484_io_data_0_in_valid = PENetwork_io_to_pes_22_in_valid; // @[pe.scala 264:34]
  assign PE_484_io_data_0_in_bits = PENetwork_io_to_pes_22_in_bits; // @[pe.scala 264:34]
  assign PE_485_clock = clock;
  assign PE_485_reset = reset;
  assign PE_485_io_data_2_sig_stat2trans = PENetwork_74_io_to_pes_1_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_485_io_data_1_in_valid = PENetwork_44_io_to_pes_1_in_valid; // @[pe.scala 264:34]
  assign PE_485_io_data_1_in_bits = PENetwork_44_io_to_pes_1_in_bits; // @[pe.scala 264:34]
  assign PE_485_io_data_0_in_valid = PENetwork_1_io_to_pes_22_in_valid; // @[pe.scala 264:34]
  assign PE_485_io_data_0_in_bits = PENetwork_1_io_to_pes_22_in_bits; // @[pe.scala 264:34]
  assign PE_486_clock = clock;
  assign PE_486_reset = reset;
  assign PE_486_io_data_2_sig_stat2trans = PENetwork_74_io_to_pes_2_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_486_io_data_1_in_valid = PENetwork_44_io_to_pes_2_in_valid; // @[pe.scala 264:34]
  assign PE_486_io_data_1_in_bits = PENetwork_44_io_to_pes_2_in_bits; // @[pe.scala 264:34]
  assign PE_486_io_data_0_in_valid = PENetwork_2_io_to_pes_22_in_valid; // @[pe.scala 264:34]
  assign PE_486_io_data_0_in_bits = PENetwork_2_io_to_pes_22_in_bits; // @[pe.scala 264:34]
  assign PE_487_clock = clock;
  assign PE_487_reset = reset;
  assign PE_487_io_data_2_sig_stat2trans = PENetwork_74_io_to_pes_3_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_487_io_data_1_in_valid = PENetwork_44_io_to_pes_3_in_valid; // @[pe.scala 264:34]
  assign PE_487_io_data_1_in_bits = PENetwork_44_io_to_pes_3_in_bits; // @[pe.scala 264:34]
  assign PE_487_io_data_0_in_valid = PENetwork_3_io_to_pes_22_in_valid; // @[pe.scala 264:34]
  assign PE_487_io_data_0_in_bits = PENetwork_3_io_to_pes_22_in_bits; // @[pe.scala 264:34]
  assign PE_488_clock = clock;
  assign PE_488_reset = reset;
  assign PE_488_io_data_2_sig_stat2trans = PENetwork_74_io_to_pes_4_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_488_io_data_1_in_valid = PENetwork_44_io_to_pes_4_in_valid; // @[pe.scala 264:34]
  assign PE_488_io_data_1_in_bits = PENetwork_44_io_to_pes_4_in_bits; // @[pe.scala 264:34]
  assign PE_488_io_data_0_in_valid = PENetwork_4_io_to_pes_22_in_valid; // @[pe.scala 264:34]
  assign PE_488_io_data_0_in_bits = PENetwork_4_io_to_pes_22_in_bits; // @[pe.scala 264:34]
  assign PE_489_clock = clock;
  assign PE_489_reset = reset;
  assign PE_489_io_data_2_sig_stat2trans = PENetwork_74_io_to_pes_5_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_489_io_data_1_in_valid = PENetwork_44_io_to_pes_5_in_valid; // @[pe.scala 264:34]
  assign PE_489_io_data_1_in_bits = PENetwork_44_io_to_pes_5_in_bits; // @[pe.scala 264:34]
  assign PE_489_io_data_0_in_valid = PENetwork_5_io_to_pes_22_in_valid; // @[pe.scala 264:34]
  assign PE_489_io_data_0_in_bits = PENetwork_5_io_to_pes_22_in_bits; // @[pe.scala 264:34]
  assign PE_490_clock = clock;
  assign PE_490_reset = reset;
  assign PE_490_io_data_2_sig_stat2trans = PENetwork_74_io_to_pes_6_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_490_io_data_1_in_valid = PENetwork_44_io_to_pes_6_in_valid; // @[pe.scala 264:34]
  assign PE_490_io_data_1_in_bits = PENetwork_44_io_to_pes_6_in_bits; // @[pe.scala 264:34]
  assign PE_490_io_data_0_in_valid = PENetwork_6_io_to_pes_22_in_valid; // @[pe.scala 264:34]
  assign PE_490_io_data_0_in_bits = PENetwork_6_io_to_pes_22_in_bits; // @[pe.scala 264:34]
  assign PE_491_clock = clock;
  assign PE_491_reset = reset;
  assign PE_491_io_data_2_sig_stat2trans = PENetwork_74_io_to_pes_7_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_491_io_data_1_in_valid = PENetwork_44_io_to_pes_7_in_valid; // @[pe.scala 264:34]
  assign PE_491_io_data_1_in_bits = PENetwork_44_io_to_pes_7_in_bits; // @[pe.scala 264:34]
  assign PE_491_io_data_0_in_valid = PENetwork_7_io_to_pes_22_in_valid; // @[pe.scala 264:34]
  assign PE_491_io_data_0_in_bits = PENetwork_7_io_to_pes_22_in_bits; // @[pe.scala 264:34]
  assign PE_492_clock = clock;
  assign PE_492_reset = reset;
  assign PE_492_io_data_2_sig_stat2trans = PENetwork_74_io_to_pes_8_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_492_io_data_1_in_valid = PENetwork_44_io_to_pes_8_in_valid; // @[pe.scala 264:34]
  assign PE_492_io_data_1_in_bits = PENetwork_44_io_to_pes_8_in_bits; // @[pe.scala 264:34]
  assign PE_492_io_data_0_in_valid = PENetwork_8_io_to_pes_22_in_valid; // @[pe.scala 264:34]
  assign PE_492_io_data_0_in_bits = PENetwork_8_io_to_pes_22_in_bits; // @[pe.scala 264:34]
  assign PE_493_clock = clock;
  assign PE_493_reset = reset;
  assign PE_493_io_data_2_sig_stat2trans = PENetwork_74_io_to_pes_9_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_493_io_data_1_in_valid = PENetwork_44_io_to_pes_9_in_valid; // @[pe.scala 264:34]
  assign PE_493_io_data_1_in_bits = PENetwork_44_io_to_pes_9_in_bits; // @[pe.scala 264:34]
  assign PE_493_io_data_0_in_valid = PENetwork_9_io_to_pes_22_in_valid; // @[pe.scala 264:34]
  assign PE_493_io_data_0_in_bits = PENetwork_9_io_to_pes_22_in_bits; // @[pe.scala 264:34]
  assign PE_494_clock = clock;
  assign PE_494_reset = reset;
  assign PE_494_io_data_2_sig_stat2trans = PENetwork_74_io_to_pes_10_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_494_io_data_1_in_valid = PENetwork_44_io_to_pes_10_in_valid; // @[pe.scala 264:34]
  assign PE_494_io_data_1_in_bits = PENetwork_44_io_to_pes_10_in_bits; // @[pe.scala 264:34]
  assign PE_494_io_data_0_in_valid = PENetwork_10_io_to_pes_22_in_valid; // @[pe.scala 264:34]
  assign PE_494_io_data_0_in_bits = PENetwork_10_io_to_pes_22_in_bits; // @[pe.scala 264:34]
  assign PE_495_clock = clock;
  assign PE_495_reset = reset;
  assign PE_495_io_data_2_sig_stat2trans = PENetwork_74_io_to_pes_11_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_495_io_data_1_in_valid = PENetwork_44_io_to_pes_11_in_valid; // @[pe.scala 264:34]
  assign PE_495_io_data_1_in_bits = PENetwork_44_io_to_pes_11_in_bits; // @[pe.scala 264:34]
  assign PE_495_io_data_0_in_valid = PENetwork_11_io_to_pes_22_in_valid; // @[pe.scala 264:34]
  assign PE_495_io_data_0_in_bits = PENetwork_11_io_to_pes_22_in_bits; // @[pe.scala 264:34]
  assign PE_496_clock = clock;
  assign PE_496_reset = reset;
  assign PE_496_io_data_2_sig_stat2trans = PENetwork_74_io_to_pes_12_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_496_io_data_1_in_valid = PENetwork_44_io_to_pes_12_in_valid; // @[pe.scala 264:34]
  assign PE_496_io_data_1_in_bits = PENetwork_44_io_to_pes_12_in_bits; // @[pe.scala 264:34]
  assign PE_496_io_data_0_in_valid = PENetwork_12_io_to_pes_22_in_valid; // @[pe.scala 264:34]
  assign PE_496_io_data_0_in_bits = PENetwork_12_io_to_pes_22_in_bits; // @[pe.scala 264:34]
  assign PE_497_clock = clock;
  assign PE_497_reset = reset;
  assign PE_497_io_data_2_sig_stat2trans = PENetwork_74_io_to_pes_13_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_497_io_data_1_in_valid = PENetwork_44_io_to_pes_13_in_valid; // @[pe.scala 264:34]
  assign PE_497_io_data_1_in_bits = PENetwork_44_io_to_pes_13_in_bits; // @[pe.scala 264:34]
  assign PE_497_io_data_0_in_valid = PENetwork_13_io_to_pes_22_in_valid; // @[pe.scala 264:34]
  assign PE_497_io_data_0_in_bits = PENetwork_13_io_to_pes_22_in_bits; // @[pe.scala 264:34]
  assign PE_498_clock = clock;
  assign PE_498_reset = reset;
  assign PE_498_io_data_2_sig_stat2trans = PENetwork_74_io_to_pes_14_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_498_io_data_1_in_valid = PENetwork_44_io_to_pes_14_in_valid; // @[pe.scala 264:34]
  assign PE_498_io_data_1_in_bits = PENetwork_44_io_to_pes_14_in_bits; // @[pe.scala 264:34]
  assign PE_498_io_data_0_in_valid = PENetwork_14_io_to_pes_22_in_valid; // @[pe.scala 264:34]
  assign PE_498_io_data_0_in_bits = PENetwork_14_io_to_pes_22_in_bits; // @[pe.scala 264:34]
  assign PE_499_clock = clock;
  assign PE_499_reset = reset;
  assign PE_499_io_data_2_sig_stat2trans = PENetwork_74_io_to_pes_15_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_499_io_data_1_in_valid = PENetwork_44_io_to_pes_15_in_valid; // @[pe.scala 264:34]
  assign PE_499_io_data_1_in_bits = PENetwork_44_io_to_pes_15_in_bits; // @[pe.scala 264:34]
  assign PE_499_io_data_0_in_valid = PENetwork_15_io_to_pes_22_in_valid; // @[pe.scala 264:34]
  assign PE_499_io_data_0_in_bits = PENetwork_15_io_to_pes_22_in_bits; // @[pe.scala 264:34]
  assign PE_500_clock = clock;
  assign PE_500_reset = reset;
  assign PE_500_io_data_2_sig_stat2trans = PENetwork_74_io_to_pes_16_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_500_io_data_1_in_valid = PENetwork_44_io_to_pes_16_in_valid; // @[pe.scala 264:34]
  assign PE_500_io_data_1_in_bits = PENetwork_44_io_to_pes_16_in_bits; // @[pe.scala 264:34]
  assign PE_500_io_data_0_in_valid = PENetwork_16_io_to_pes_22_in_valid; // @[pe.scala 264:34]
  assign PE_500_io_data_0_in_bits = PENetwork_16_io_to_pes_22_in_bits; // @[pe.scala 264:34]
  assign PE_501_clock = clock;
  assign PE_501_reset = reset;
  assign PE_501_io_data_2_sig_stat2trans = PENetwork_74_io_to_pes_17_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_501_io_data_1_in_valid = PENetwork_44_io_to_pes_17_in_valid; // @[pe.scala 264:34]
  assign PE_501_io_data_1_in_bits = PENetwork_44_io_to_pes_17_in_bits; // @[pe.scala 264:34]
  assign PE_501_io_data_0_in_valid = PENetwork_17_io_to_pes_22_in_valid; // @[pe.scala 264:34]
  assign PE_501_io_data_0_in_bits = PENetwork_17_io_to_pes_22_in_bits; // @[pe.scala 264:34]
  assign PE_502_clock = clock;
  assign PE_502_reset = reset;
  assign PE_502_io_data_2_sig_stat2trans = PENetwork_74_io_to_pes_18_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_502_io_data_1_in_valid = PENetwork_44_io_to_pes_18_in_valid; // @[pe.scala 264:34]
  assign PE_502_io_data_1_in_bits = PENetwork_44_io_to_pes_18_in_bits; // @[pe.scala 264:34]
  assign PE_502_io_data_0_in_valid = PENetwork_18_io_to_pes_22_in_valid; // @[pe.scala 264:34]
  assign PE_502_io_data_0_in_bits = PENetwork_18_io_to_pes_22_in_bits; // @[pe.scala 264:34]
  assign PE_503_clock = clock;
  assign PE_503_reset = reset;
  assign PE_503_io_data_2_sig_stat2trans = PENetwork_74_io_to_pes_19_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_503_io_data_1_in_valid = PENetwork_44_io_to_pes_19_in_valid; // @[pe.scala 264:34]
  assign PE_503_io_data_1_in_bits = PENetwork_44_io_to_pes_19_in_bits; // @[pe.scala 264:34]
  assign PE_503_io_data_0_in_valid = PENetwork_19_io_to_pes_22_in_valid; // @[pe.scala 264:34]
  assign PE_503_io_data_0_in_bits = PENetwork_19_io_to_pes_22_in_bits; // @[pe.scala 264:34]
  assign PE_504_clock = clock;
  assign PE_504_reset = reset;
  assign PE_504_io_data_2_sig_stat2trans = PENetwork_74_io_to_pes_20_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_504_io_data_1_in_valid = PENetwork_44_io_to_pes_20_in_valid; // @[pe.scala 264:34]
  assign PE_504_io_data_1_in_bits = PENetwork_44_io_to_pes_20_in_bits; // @[pe.scala 264:34]
  assign PE_504_io_data_0_in_valid = PENetwork_20_io_to_pes_22_in_valid; // @[pe.scala 264:34]
  assign PE_504_io_data_0_in_bits = PENetwork_20_io_to_pes_22_in_bits; // @[pe.scala 264:34]
  assign PE_505_clock = clock;
  assign PE_505_reset = reset;
  assign PE_505_io_data_2_sig_stat2trans = PENetwork_74_io_to_pes_21_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_505_io_data_1_in_valid = PENetwork_44_io_to_pes_21_in_valid; // @[pe.scala 264:34]
  assign PE_505_io_data_1_in_bits = PENetwork_44_io_to_pes_21_in_bits; // @[pe.scala 264:34]
  assign PE_505_io_data_0_in_valid = PENetwork_21_io_to_pes_22_in_valid; // @[pe.scala 264:34]
  assign PE_505_io_data_0_in_bits = PENetwork_21_io_to_pes_22_in_bits; // @[pe.scala 264:34]
  assign PE_506_clock = clock;
  assign PE_506_reset = reset;
  assign PE_506_io_data_2_sig_stat2trans = PENetwork_75_io_to_pes_0_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_506_io_data_1_in_valid = PENetwork_45_io_to_pes_0_in_valid; // @[pe.scala 264:34]
  assign PE_506_io_data_1_in_bits = PENetwork_45_io_to_pes_0_in_bits; // @[pe.scala 264:34]
  assign PE_506_io_data_0_in_valid = PENetwork_io_to_pes_23_in_valid; // @[pe.scala 264:34]
  assign PE_506_io_data_0_in_bits = PENetwork_io_to_pes_23_in_bits; // @[pe.scala 264:34]
  assign PE_507_clock = clock;
  assign PE_507_reset = reset;
  assign PE_507_io_data_2_sig_stat2trans = PENetwork_75_io_to_pes_1_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_507_io_data_1_in_valid = PENetwork_45_io_to_pes_1_in_valid; // @[pe.scala 264:34]
  assign PE_507_io_data_1_in_bits = PENetwork_45_io_to_pes_1_in_bits; // @[pe.scala 264:34]
  assign PE_507_io_data_0_in_valid = PENetwork_1_io_to_pes_23_in_valid; // @[pe.scala 264:34]
  assign PE_507_io_data_0_in_bits = PENetwork_1_io_to_pes_23_in_bits; // @[pe.scala 264:34]
  assign PE_508_clock = clock;
  assign PE_508_reset = reset;
  assign PE_508_io_data_2_sig_stat2trans = PENetwork_75_io_to_pes_2_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_508_io_data_1_in_valid = PENetwork_45_io_to_pes_2_in_valid; // @[pe.scala 264:34]
  assign PE_508_io_data_1_in_bits = PENetwork_45_io_to_pes_2_in_bits; // @[pe.scala 264:34]
  assign PE_508_io_data_0_in_valid = PENetwork_2_io_to_pes_23_in_valid; // @[pe.scala 264:34]
  assign PE_508_io_data_0_in_bits = PENetwork_2_io_to_pes_23_in_bits; // @[pe.scala 264:34]
  assign PE_509_clock = clock;
  assign PE_509_reset = reset;
  assign PE_509_io_data_2_sig_stat2trans = PENetwork_75_io_to_pes_3_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_509_io_data_1_in_valid = PENetwork_45_io_to_pes_3_in_valid; // @[pe.scala 264:34]
  assign PE_509_io_data_1_in_bits = PENetwork_45_io_to_pes_3_in_bits; // @[pe.scala 264:34]
  assign PE_509_io_data_0_in_valid = PENetwork_3_io_to_pes_23_in_valid; // @[pe.scala 264:34]
  assign PE_509_io_data_0_in_bits = PENetwork_3_io_to_pes_23_in_bits; // @[pe.scala 264:34]
  assign PE_510_clock = clock;
  assign PE_510_reset = reset;
  assign PE_510_io_data_2_sig_stat2trans = PENetwork_75_io_to_pes_4_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_510_io_data_1_in_valid = PENetwork_45_io_to_pes_4_in_valid; // @[pe.scala 264:34]
  assign PE_510_io_data_1_in_bits = PENetwork_45_io_to_pes_4_in_bits; // @[pe.scala 264:34]
  assign PE_510_io_data_0_in_valid = PENetwork_4_io_to_pes_23_in_valid; // @[pe.scala 264:34]
  assign PE_510_io_data_0_in_bits = PENetwork_4_io_to_pes_23_in_bits; // @[pe.scala 264:34]
  assign PE_511_clock = clock;
  assign PE_511_reset = reset;
  assign PE_511_io_data_2_sig_stat2trans = PENetwork_75_io_to_pes_5_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_511_io_data_1_in_valid = PENetwork_45_io_to_pes_5_in_valid; // @[pe.scala 264:34]
  assign PE_511_io_data_1_in_bits = PENetwork_45_io_to_pes_5_in_bits; // @[pe.scala 264:34]
  assign PE_511_io_data_0_in_valid = PENetwork_5_io_to_pes_23_in_valid; // @[pe.scala 264:34]
  assign PE_511_io_data_0_in_bits = PENetwork_5_io_to_pes_23_in_bits; // @[pe.scala 264:34]
  assign PE_512_clock = clock;
  assign PE_512_reset = reset;
  assign PE_512_io_data_2_sig_stat2trans = PENetwork_75_io_to_pes_6_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_512_io_data_1_in_valid = PENetwork_45_io_to_pes_6_in_valid; // @[pe.scala 264:34]
  assign PE_512_io_data_1_in_bits = PENetwork_45_io_to_pes_6_in_bits; // @[pe.scala 264:34]
  assign PE_512_io_data_0_in_valid = PENetwork_6_io_to_pes_23_in_valid; // @[pe.scala 264:34]
  assign PE_512_io_data_0_in_bits = PENetwork_6_io_to_pes_23_in_bits; // @[pe.scala 264:34]
  assign PE_513_clock = clock;
  assign PE_513_reset = reset;
  assign PE_513_io_data_2_sig_stat2trans = PENetwork_75_io_to_pes_7_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_513_io_data_1_in_valid = PENetwork_45_io_to_pes_7_in_valid; // @[pe.scala 264:34]
  assign PE_513_io_data_1_in_bits = PENetwork_45_io_to_pes_7_in_bits; // @[pe.scala 264:34]
  assign PE_513_io_data_0_in_valid = PENetwork_7_io_to_pes_23_in_valid; // @[pe.scala 264:34]
  assign PE_513_io_data_0_in_bits = PENetwork_7_io_to_pes_23_in_bits; // @[pe.scala 264:34]
  assign PE_514_clock = clock;
  assign PE_514_reset = reset;
  assign PE_514_io_data_2_sig_stat2trans = PENetwork_75_io_to_pes_8_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_514_io_data_1_in_valid = PENetwork_45_io_to_pes_8_in_valid; // @[pe.scala 264:34]
  assign PE_514_io_data_1_in_bits = PENetwork_45_io_to_pes_8_in_bits; // @[pe.scala 264:34]
  assign PE_514_io_data_0_in_valid = PENetwork_8_io_to_pes_23_in_valid; // @[pe.scala 264:34]
  assign PE_514_io_data_0_in_bits = PENetwork_8_io_to_pes_23_in_bits; // @[pe.scala 264:34]
  assign PE_515_clock = clock;
  assign PE_515_reset = reset;
  assign PE_515_io_data_2_sig_stat2trans = PENetwork_75_io_to_pes_9_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_515_io_data_1_in_valid = PENetwork_45_io_to_pes_9_in_valid; // @[pe.scala 264:34]
  assign PE_515_io_data_1_in_bits = PENetwork_45_io_to_pes_9_in_bits; // @[pe.scala 264:34]
  assign PE_515_io_data_0_in_valid = PENetwork_9_io_to_pes_23_in_valid; // @[pe.scala 264:34]
  assign PE_515_io_data_0_in_bits = PENetwork_9_io_to_pes_23_in_bits; // @[pe.scala 264:34]
  assign PE_516_clock = clock;
  assign PE_516_reset = reset;
  assign PE_516_io_data_2_sig_stat2trans = PENetwork_75_io_to_pes_10_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_516_io_data_1_in_valid = PENetwork_45_io_to_pes_10_in_valid; // @[pe.scala 264:34]
  assign PE_516_io_data_1_in_bits = PENetwork_45_io_to_pes_10_in_bits; // @[pe.scala 264:34]
  assign PE_516_io_data_0_in_valid = PENetwork_10_io_to_pes_23_in_valid; // @[pe.scala 264:34]
  assign PE_516_io_data_0_in_bits = PENetwork_10_io_to_pes_23_in_bits; // @[pe.scala 264:34]
  assign PE_517_clock = clock;
  assign PE_517_reset = reset;
  assign PE_517_io_data_2_sig_stat2trans = PENetwork_75_io_to_pes_11_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_517_io_data_1_in_valid = PENetwork_45_io_to_pes_11_in_valid; // @[pe.scala 264:34]
  assign PE_517_io_data_1_in_bits = PENetwork_45_io_to_pes_11_in_bits; // @[pe.scala 264:34]
  assign PE_517_io_data_0_in_valid = PENetwork_11_io_to_pes_23_in_valid; // @[pe.scala 264:34]
  assign PE_517_io_data_0_in_bits = PENetwork_11_io_to_pes_23_in_bits; // @[pe.scala 264:34]
  assign PE_518_clock = clock;
  assign PE_518_reset = reset;
  assign PE_518_io_data_2_sig_stat2trans = PENetwork_75_io_to_pes_12_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_518_io_data_1_in_valid = PENetwork_45_io_to_pes_12_in_valid; // @[pe.scala 264:34]
  assign PE_518_io_data_1_in_bits = PENetwork_45_io_to_pes_12_in_bits; // @[pe.scala 264:34]
  assign PE_518_io_data_0_in_valid = PENetwork_12_io_to_pes_23_in_valid; // @[pe.scala 264:34]
  assign PE_518_io_data_0_in_bits = PENetwork_12_io_to_pes_23_in_bits; // @[pe.scala 264:34]
  assign PE_519_clock = clock;
  assign PE_519_reset = reset;
  assign PE_519_io_data_2_sig_stat2trans = PENetwork_75_io_to_pes_13_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_519_io_data_1_in_valid = PENetwork_45_io_to_pes_13_in_valid; // @[pe.scala 264:34]
  assign PE_519_io_data_1_in_bits = PENetwork_45_io_to_pes_13_in_bits; // @[pe.scala 264:34]
  assign PE_519_io_data_0_in_valid = PENetwork_13_io_to_pes_23_in_valid; // @[pe.scala 264:34]
  assign PE_519_io_data_0_in_bits = PENetwork_13_io_to_pes_23_in_bits; // @[pe.scala 264:34]
  assign PE_520_clock = clock;
  assign PE_520_reset = reset;
  assign PE_520_io_data_2_sig_stat2trans = PENetwork_75_io_to_pes_14_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_520_io_data_1_in_valid = PENetwork_45_io_to_pes_14_in_valid; // @[pe.scala 264:34]
  assign PE_520_io_data_1_in_bits = PENetwork_45_io_to_pes_14_in_bits; // @[pe.scala 264:34]
  assign PE_520_io_data_0_in_valid = PENetwork_14_io_to_pes_23_in_valid; // @[pe.scala 264:34]
  assign PE_520_io_data_0_in_bits = PENetwork_14_io_to_pes_23_in_bits; // @[pe.scala 264:34]
  assign PE_521_clock = clock;
  assign PE_521_reset = reset;
  assign PE_521_io_data_2_sig_stat2trans = PENetwork_75_io_to_pes_15_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_521_io_data_1_in_valid = PENetwork_45_io_to_pes_15_in_valid; // @[pe.scala 264:34]
  assign PE_521_io_data_1_in_bits = PENetwork_45_io_to_pes_15_in_bits; // @[pe.scala 264:34]
  assign PE_521_io_data_0_in_valid = PENetwork_15_io_to_pes_23_in_valid; // @[pe.scala 264:34]
  assign PE_521_io_data_0_in_bits = PENetwork_15_io_to_pes_23_in_bits; // @[pe.scala 264:34]
  assign PE_522_clock = clock;
  assign PE_522_reset = reset;
  assign PE_522_io_data_2_sig_stat2trans = PENetwork_75_io_to_pes_16_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_522_io_data_1_in_valid = PENetwork_45_io_to_pes_16_in_valid; // @[pe.scala 264:34]
  assign PE_522_io_data_1_in_bits = PENetwork_45_io_to_pes_16_in_bits; // @[pe.scala 264:34]
  assign PE_522_io_data_0_in_valid = PENetwork_16_io_to_pes_23_in_valid; // @[pe.scala 264:34]
  assign PE_522_io_data_0_in_bits = PENetwork_16_io_to_pes_23_in_bits; // @[pe.scala 264:34]
  assign PE_523_clock = clock;
  assign PE_523_reset = reset;
  assign PE_523_io_data_2_sig_stat2trans = PENetwork_75_io_to_pes_17_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_523_io_data_1_in_valid = PENetwork_45_io_to_pes_17_in_valid; // @[pe.scala 264:34]
  assign PE_523_io_data_1_in_bits = PENetwork_45_io_to_pes_17_in_bits; // @[pe.scala 264:34]
  assign PE_523_io_data_0_in_valid = PENetwork_17_io_to_pes_23_in_valid; // @[pe.scala 264:34]
  assign PE_523_io_data_0_in_bits = PENetwork_17_io_to_pes_23_in_bits; // @[pe.scala 264:34]
  assign PE_524_clock = clock;
  assign PE_524_reset = reset;
  assign PE_524_io_data_2_sig_stat2trans = PENetwork_75_io_to_pes_18_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_524_io_data_1_in_valid = PENetwork_45_io_to_pes_18_in_valid; // @[pe.scala 264:34]
  assign PE_524_io_data_1_in_bits = PENetwork_45_io_to_pes_18_in_bits; // @[pe.scala 264:34]
  assign PE_524_io_data_0_in_valid = PENetwork_18_io_to_pes_23_in_valid; // @[pe.scala 264:34]
  assign PE_524_io_data_0_in_bits = PENetwork_18_io_to_pes_23_in_bits; // @[pe.scala 264:34]
  assign PE_525_clock = clock;
  assign PE_525_reset = reset;
  assign PE_525_io_data_2_sig_stat2trans = PENetwork_75_io_to_pes_19_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_525_io_data_1_in_valid = PENetwork_45_io_to_pes_19_in_valid; // @[pe.scala 264:34]
  assign PE_525_io_data_1_in_bits = PENetwork_45_io_to_pes_19_in_bits; // @[pe.scala 264:34]
  assign PE_525_io_data_0_in_valid = PENetwork_19_io_to_pes_23_in_valid; // @[pe.scala 264:34]
  assign PE_525_io_data_0_in_bits = PENetwork_19_io_to_pes_23_in_bits; // @[pe.scala 264:34]
  assign PE_526_clock = clock;
  assign PE_526_reset = reset;
  assign PE_526_io_data_2_sig_stat2trans = PENetwork_75_io_to_pes_20_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_526_io_data_1_in_valid = PENetwork_45_io_to_pes_20_in_valid; // @[pe.scala 264:34]
  assign PE_526_io_data_1_in_bits = PENetwork_45_io_to_pes_20_in_bits; // @[pe.scala 264:34]
  assign PE_526_io_data_0_in_valid = PENetwork_20_io_to_pes_23_in_valid; // @[pe.scala 264:34]
  assign PE_526_io_data_0_in_bits = PENetwork_20_io_to_pes_23_in_bits; // @[pe.scala 264:34]
  assign PE_527_clock = clock;
  assign PE_527_reset = reset;
  assign PE_527_io_data_2_sig_stat2trans = PENetwork_75_io_to_pes_21_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_527_io_data_1_in_valid = PENetwork_45_io_to_pes_21_in_valid; // @[pe.scala 264:34]
  assign PE_527_io_data_1_in_bits = PENetwork_45_io_to_pes_21_in_bits; // @[pe.scala 264:34]
  assign PE_527_io_data_0_in_valid = PENetwork_21_io_to_pes_23_in_valid; // @[pe.scala 264:34]
  assign PE_527_io_data_0_in_bits = PENetwork_21_io_to_pes_23_in_bits; // @[pe.scala 264:34]
  assign PE_528_clock = clock;
  assign PE_528_reset = reset;
  assign PE_528_io_data_2_sig_stat2trans = PENetwork_76_io_to_pes_0_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_528_io_data_1_in_valid = PENetwork_46_io_to_pes_0_in_valid; // @[pe.scala 264:34]
  assign PE_528_io_data_1_in_bits = PENetwork_46_io_to_pes_0_in_bits; // @[pe.scala 264:34]
  assign PE_528_io_data_0_in_valid = PENetwork_io_to_pes_24_in_valid; // @[pe.scala 264:34]
  assign PE_528_io_data_0_in_bits = PENetwork_io_to_pes_24_in_bits; // @[pe.scala 264:34]
  assign PE_529_clock = clock;
  assign PE_529_reset = reset;
  assign PE_529_io_data_2_sig_stat2trans = PENetwork_76_io_to_pes_1_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_529_io_data_1_in_valid = PENetwork_46_io_to_pes_1_in_valid; // @[pe.scala 264:34]
  assign PE_529_io_data_1_in_bits = PENetwork_46_io_to_pes_1_in_bits; // @[pe.scala 264:34]
  assign PE_529_io_data_0_in_valid = PENetwork_1_io_to_pes_24_in_valid; // @[pe.scala 264:34]
  assign PE_529_io_data_0_in_bits = PENetwork_1_io_to_pes_24_in_bits; // @[pe.scala 264:34]
  assign PE_530_clock = clock;
  assign PE_530_reset = reset;
  assign PE_530_io_data_2_sig_stat2trans = PENetwork_76_io_to_pes_2_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_530_io_data_1_in_valid = PENetwork_46_io_to_pes_2_in_valid; // @[pe.scala 264:34]
  assign PE_530_io_data_1_in_bits = PENetwork_46_io_to_pes_2_in_bits; // @[pe.scala 264:34]
  assign PE_530_io_data_0_in_valid = PENetwork_2_io_to_pes_24_in_valid; // @[pe.scala 264:34]
  assign PE_530_io_data_0_in_bits = PENetwork_2_io_to_pes_24_in_bits; // @[pe.scala 264:34]
  assign PE_531_clock = clock;
  assign PE_531_reset = reset;
  assign PE_531_io_data_2_sig_stat2trans = PENetwork_76_io_to_pes_3_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_531_io_data_1_in_valid = PENetwork_46_io_to_pes_3_in_valid; // @[pe.scala 264:34]
  assign PE_531_io_data_1_in_bits = PENetwork_46_io_to_pes_3_in_bits; // @[pe.scala 264:34]
  assign PE_531_io_data_0_in_valid = PENetwork_3_io_to_pes_24_in_valid; // @[pe.scala 264:34]
  assign PE_531_io_data_0_in_bits = PENetwork_3_io_to_pes_24_in_bits; // @[pe.scala 264:34]
  assign PE_532_clock = clock;
  assign PE_532_reset = reset;
  assign PE_532_io_data_2_sig_stat2trans = PENetwork_76_io_to_pes_4_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_532_io_data_1_in_valid = PENetwork_46_io_to_pes_4_in_valid; // @[pe.scala 264:34]
  assign PE_532_io_data_1_in_bits = PENetwork_46_io_to_pes_4_in_bits; // @[pe.scala 264:34]
  assign PE_532_io_data_0_in_valid = PENetwork_4_io_to_pes_24_in_valid; // @[pe.scala 264:34]
  assign PE_532_io_data_0_in_bits = PENetwork_4_io_to_pes_24_in_bits; // @[pe.scala 264:34]
  assign PE_533_clock = clock;
  assign PE_533_reset = reset;
  assign PE_533_io_data_2_sig_stat2trans = PENetwork_76_io_to_pes_5_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_533_io_data_1_in_valid = PENetwork_46_io_to_pes_5_in_valid; // @[pe.scala 264:34]
  assign PE_533_io_data_1_in_bits = PENetwork_46_io_to_pes_5_in_bits; // @[pe.scala 264:34]
  assign PE_533_io_data_0_in_valid = PENetwork_5_io_to_pes_24_in_valid; // @[pe.scala 264:34]
  assign PE_533_io_data_0_in_bits = PENetwork_5_io_to_pes_24_in_bits; // @[pe.scala 264:34]
  assign PE_534_clock = clock;
  assign PE_534_reset = reset;
  assign PE_534_io_data_2_sig_stat2trans = PENetwork_76_io_to_pes_6_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_534_io_data_1_in_valid = PENetwork_46_io_to_pes_6_in_valid; // @[pe.scala 264:34]
  assign PE_534_io_data_1_in_bits = PENetwork_46_io_to_pes_6_in_bits; // @[pe.scala 264:34]
  assign PE_534_io_data_0_in_valid = PENetwork_6_io_to_pes_24_in_valid; // @[pe.scala 264:34]
  assign PE_534_io_data_0_in_bits = PENetwork_6_io_to_pes_24_in_bits; // @[pe.scala 264:34]
  assign PE_535_clock = clock;
  assign PE_535_reset = reset;
  assign PE_535_io_data_2_sig_stat2trans = PENetwork_76_io_to_pes_7_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_535_io_data_1_in_valid = PENetwork_46_io_to_pes_7_in_valid; // @[pe.scala 264:34]
  assign PE_535_io_data_1_in_bits = PENetwork_46_io_to_pes_7_in_bits; // @[pe.scala 264:34]
  assign PE_535_io_data_0_in_valid = PENetwork_7_io_to_pes_24_in_valid; // @[pe.scala 264:34]
  assign PE_535_io_data_0_in_bits = PENetwork_7_io_to_pes_24_in_bits; // @[pe.scala 264:34]
  assign PE_536_clock = clock;
  assign PE_536_reset = reset;
  assign PE_536_io_data_2_sig_stat2trans = PENetwork_76_io_to_pes_8_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_536_io_data_1_in_valid = PENetwork_46_io_to_pes_8_in_valid; // @[pe.scala 264:34]
  assign PE_536_io_data_1_in_bits = PENetwork_46_io_to_pes_8_in_bits; // @[pe.scala 264:34]
  assign PE_536_io_data_0_in_valid = PENetwork_8_io_to_pes_24_in_valid; // @[pe.scala 264:34]
  assign PE_536_io_data_0_in_bits = PENetwork_8_io_to_pes_24_in_bits; // @[pe.scala 264:34]
  assign PE_537_clock = clock;
  assign PE_537_reset = reset;
  assign PE_537_io_data_2_sig_stat2trans = PENetwork_76_io_to_pes_9_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_537_io_data_1_in_valid = PENetwork_46_io_to_pes_9_in_valid; // @[pe.scala 264:34]
  assign PE_537_io_data_1_in_bits = PENetwork_46_io_to_pes_9_in_bits; // @[pe.scala 264:34]
  assign PE_537_io_data_0_in_valid = PENetwork_9_io_to_pes_24_in_valid; // @[pe.scala 264:34]
  assign PE_537_io_data_0_in_bits = PENetwork_9_io_to_pes_24_in_bits; // @[pe.scala 264:34]
  assign PE_538_clock = clock;
  assign PE_538_reset = reset;
  assign PE_538_io_data_2_sig_stat2trans = PENetwork_76_io_to_pes_10_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_538_io_data_1_in_valid = PENetwork_46_io_to_pes_10_in_valid; // @[pe.scala 264:34]
  assign PE_538_io_data_1_in_bits = PENetwork_46_io_to_pes_10_in_bits; // @[pe.scala 264:34]
  assign PE_538_io_data_0_in_valid = PENetwork_10_io_to_pes_24_in_valid; // @[pe.scala 264:34]
  assign PE_538_io_data_0_in_bits = PENetwork_10_io_to_pes_24_in_bits; // @[pe.scala 264:34]
  assign PE_539_clock = clock;
  assign PE_539_reset = reset;
  assign PE_539_io_data_2_sig_stat2trans = PENetwork_76_io_to_pes_11_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_539_io_data_1_in_valid = PENetwork_46_io_to_pes_11_in_valid; // @[pe.scala 264:34]
  assign PE_539_io_data_1_in_bits = PENetwork_46_io_to_pes_11_in_bits; // @[pe.scala 264:34]
  assign PE_539_io_data_0_in_valid = PENetwork_11_io_to_pes_24_in_valid; // @[pe.scala 264:34]
  assign PE_539_io_data_0_in_bits = PENetwork_11_io_to_pes_24_in_bits; // @[pe.scala 264:34]
  assign PE_540_clock = clock;
  assign PE_540_reset = reset;
  assign PE_540_io_data_2_sig_stat2trans = PENetwork_76_io_to_pes_12_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_540_io_data_1_in_valid = PENetwork_46_io_to_pes_12_in_valid; // @[pe.scala 264:34]
  assign PE_540_io_data_1_in_bits = PENetwork_46_io_to_pes_12_in_bits; // @[pe.scala 264:34]
  assign PE_540_io_data_0_in_valid = PENetwork_12_io_to_pes_24_in_valid; // @[pe.scala 264:34]
  assign PE_540_io_data_0_in_bits = PENetwork_12_io_to_pes_24_in_bits; // @[pe.scala 264:34]
  assign PE_541_clock = clock;
  assign PE_541_reset = reset;
  assign PE_541_io_data_2_sig_stat2trans = PENetwork_76_io_to_pes_13_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_541_io_data_1_in_valid = PENetwork_46_io_to_pes_13_in_valid; // @[pe.scala 264:34]
  assign PE_541_io_data_1_in_bits = PENetwork_46_io_to_pes_13_in_bits; // @[pe.scala 264:34]
  assign PE_541_io_data_0_in_valid = PENetwork_13_io_to_pes_24_in_valid; // @[pe.scala 264:34]
  assign PE_541_io_data_0_in_bits = PENetwork_13_io_to_pes_24_in_bits; // @[pe.scala 264:34]
  assign PE_542_clock = clock;
  assign PE_542_reset = reset;
  assign PE_542_io_data_2_sig_stat2trans = PENetwork_76_io_to_pes_14_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_542_io_data_1_in_valid = PENetwork_46_io_to_pes_14_in_valid; // @[pe.scala 264:34]
  assign PE_542_io_data_1_in_bits = PENetwork_46_io_to_pes_14_in_bits; // @[pe.scala 264:34]
  assign PE_542_io_data_0_in_valid = PENetwork_14_io_to_pes_24_in_valid; // @[pe.scala 264:34]
  assign PE_542_io_data_0_in_bits = PENetwork_14_io_to_pes_24_in_bits; // @[pe.scala 264:34]
  assign PE_543_clock = clock;
  assign PE_543_reset = reset;
  assign PE_543_io_data_2_sig_stat2trans = PENetwork_76_io_to_pes_15_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_543_io_data_1_in_valid = PENetwork_46_io_to_pes_15_in_valid; // @[pe.scala 264:34]
  assign PE_543_io_data_1_in_bits = PENetwork_46_io_to_pes_15_in_bits; // @[pe.scala 264:34]
  assign PE_543_io_data_0_in_valid = PENetwork_15_io_to_pes_24_in_valid; // @[pe.scala 264:34]
  assign PE_543_io_data_0_in_bits = PENetwork_15_io_to_pes_24_in_bits; // @[pe.scala 264:34]
  assign PE_544_clock = clock;
  assign PE_544_reset = reset;
  assign PE_544_io_data_2_sig_stat2trans = PENetwork_76_io_to_pes_16_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_544_io_data_1_in_valid = PENetwork_46_io_to_pes_16_in_valid; // @[pe.scala 264:34]
  assign PE_544_io_data_1_in_bits = PENetwork_46_io_to_pes_16_in_bits; // @[pe.scala 264:34]
  assign PE_544_io_data_0_in_valid = PENetwork_16_io_to_pes_24_in_valid; // @[pe.scala 264:34]
  assign PE_544_io_data_0_in_bits = PENetwork_16_io_to_pes_24_in_bits; // @[pe.scala 264:34]
  assign PE_545_clock = clock;
  assign PE_545_reset = reset;
  assign PE_545_io_data_2_sig_stat2trans = PENetwork_76_io_to_pes_17_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_545_io_data_1_in_valid = PENetwork_46_io_to_pes_17_in_valid; // @[pe.scala 264:34]
  assign PE_545_io_data_1_in_bits = PENetwork_46_io_to_pes_17_in_bits; // @[pe.scala 264:34]
  assign PE_545_io_data_0_in_valid = PENetwork_17_io_to_pes_24_in_valid; // @[pe.scala 264:34]
  assign PE_545_io_data_0_in_bits = PENetwork_17_io_to_pes_24_in_bits; // @[pe.scala 264:34]
  assign PE_546_clock = clock;
  assign PE_546_reset = reset;
  assign PE_546_io_data_2_sig_stat2trans = PENetwork_76_io_to_pes_18_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_546_io_data_1_in_valid = PENetwork_46_io_to_pes_18_in_valid; // @[pe.scala 264:34]
  assign PE_546_io_data_1_in_bits = PENetwork_46_io_to_pes_18_in_bits; // @[pe.scala 264:34]
  assign PE_546_io_data_0_in_valid = PENetwork_18_io_to_pes_24_in_valid; // @[pe.scala 264:34]
  assign PE_546_io_data_0_in_bits = PENetwork_18_io_to_pes_24_in_bits; // @[pe.scala 264:34]
  assign PE_547_clock = clock;
  assign PE_547_reset = reset;
  assign PE_547_io_data_2_sig_stat2trans = PENetwork_76_io_to_pes_19_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_547_io_data_1_in_valid = PENetwork_46_io_to_pes_19_in_valid; // @[pe.scala 264:34]
  assign PE_547_io_data_1_in_bits = PENetwork_46_io_to_pes_19_in_bits; // @[pe.scala 264:34]
  assign PE_547_io_data_0_in_valid = PENetwork_19_io_to_pes_24_in_valid; // @[pe.scala 264:34]
  assign PE_547_io_data_0_in_bits = PENetwork_19_io_to_pes_24_in_bits; // @[pe.scala 264:34]
  assign PE_548_clock = clock;
  assign PE_548_reset = reset;
  assign PE_548_io_data_2_sig_stat2trans = PENetwork_76_io_to_pes_20_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_548_io_data_1_in_valid = PENetwork_46_io_to_pes_20_in_valid; // @[pe.scala 264:34]
  assign PE_548_io_data_1_in_bits = PENetwork_46_io_to_pes_20_in_bits; // @[pe.scala 264:34]
  assign PE_548_io_data_0_in_valid = PENetwork_20_io_to_pes_24_in_valid; // @[pe.scala 264:34]
  assign PE_548_io_data_0_in_bits = PENetwork_20_io_to_pes_24_in_bits; // @[pe.scala 264:34]
  assign PE_549_clock = clock;
  assign PE_549_reset = reset;
  assign PE_549_io_data_2_sig_stat2trans = PENetwork_76_io_to_pes_21_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_549_io_data_1_in_valid = PENetwork_46_io_to_pes_21_in_valid; // @[pe.scala 264:34]
  assign PE_549_io_data_1_in_bits = PENetwork_46_io_to_pes_21_in_bits; // @[pe.scala 264:34]
  assign PE_549_io_data_0_in_valid = PENetwork_21_io_to_pes_24_in_valid; // @[pe.scala 264:34]
  assign PE_549_io_data_0_in_bits = PENetwork_21_io_to_pes_24_in_bits; // @[pe.scala 264:34]
  assign PE_550_clock = clock;
  assign PE_550_reset = reset;
  assign PE_550_io_data_2_sig_stat2trans = PENetwork_77_io_to_pes_0_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_550_io_data_1_in_valid = PENetwork_47_io_to_pes_0_in_valid; // @[pe.scala 264:34]
  assign PE_550_io_data_1_in_bits = PENetwork_47_io_to_pes_0_in_bits; // @[pe.scala 264:34]
  assign PE_550_io_data_0_in_valid = PENetwork_io_to_pes_25_in_valid; // @[pe.scala 264:34]
  assign PE_550_io_data_0_in_bits = PENetwork_io_to_pes_25_in_bits; // @[pe.scala 264:34]
  assign PE_551_clock = clock;
  assign PE_551_reset = reset;
  assign PE_551_io_data_2_sig_stat2trans = PENetwork_77_io_to_pes_1_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_551_io_data_1_in_valid = PENetwork_47_io_to_pes_1_in_valid; // @[pe.scala 264:34]
  assign PE_551_io_data_1_in_bits = PENetwork_47_io_to_pes_1_in_bits; // @[pe.scala 264:34]
  assign PE_551_io_data_0_in_valid = PENetwork_1_io_to_pes_25_in_valid; // @[pe.scala 264:34]
  assign PE_551_io_data_0_in_bits = PENetwork_1_io_to_pes_25_in_bits; // @[pe.scala 264:34]
  assign PE_552_clock = clock;
  assign PE_552_reset = reset;
  assign PE_552_io_data_2_sig_stat2trans = PENetwork_77_io_to_pes_2_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_552_io_data_1_in_valid = PENetwork_47_io_to_pes_2_in_valid; // @[pe.scala 264:34]
  assign PE_552_io_data_1_in_bits = PENetwork_47_io_to_pes_2_in_bits; // @[pe.scala 264:34]
  assign PE_552_io_data_0_in_valid = PENetwork_2_io_to_pes_25_in_valid; // @[pe.scala 264:34]
  assign PE_552_io_data_0_in_bits = PENetwork_2_io_to_pes_25_in_bits; // @[pe.scala 264:34]
  assign PE_553_clock = clock;
  assign PE_553_reset = reset;
  assign PE_553_io_data_2_sig_stat2trans = PENetwork_77_io_to_pes_3_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_553_io_data_1_in_valid = PENetwork_47_io_to_pes_3_in_valid; // @[pe.scala 264:34]
  assign PE_553_io_data_1_in_bits = PENetwork_47_io_to_pes_3_in_bits; // @[pe.scala 264:34]
  assign PE_553_io_data_0_in_valid = PENetwork_3_io_to_pes_25_in_valid; // @[pe.scala 264:34]
  assign PE_553_io_data_0_in_bits = PENetwork_3_io_to_pes_25_in_bits; // @[pe.scala 264:34]
  assign PE_554_clock = clock;
  assign PE_554_reset = reset;
  assign PE_554_io_data_2_sig_stat2trans = PENetwork_77_io_to_pes_4_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_554_io_data_1_in_valid = PENetwork_47_io_to_pes_4_in_valid; // @[pe.scala 264:34]
  assign PE_554_io_data_1_in_bits = PENetwork_47_io_to_pes_4_in_bits; // @[pe.scala 264:34]
  assign PE_554_io_data_0_in_valid = PENetwork_4_io_to_pes_25_in_valid; // @[pe.scala 264:34]
  assign PE_554_io_data_0_in_bits = PENetwork_4_io_to_pes_25_in_bits; // @[pe.scala 264:34]
  assign PE_555_clock = clock;
  assign PE_555_reset = reset;
  assign PE_555_io_data_2_sig_stat2trans = PENetwork_77_io_to_pes_5_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_555_io_data_1_in_valid = PENetwork_47_io_to_pes_5_in_valid; // @[pe.scala 264:34]
  assign PE_555_io_data_1_in_bits = PENetwork_47_io_to_pes_5_in_bits; // @[pe.scala 264:34]
  assign PE_555_io_data_0_in_valid = PENetwork_5_io_to_pes_25_in_valid; // @[pe.scala 264:34]
  assign PE_555_io_data_0_in_bits = PENetwork_5_io_to_pes_25_in_bits; // @[pe.scala 264:34]
  assign PE_556_clock = clock;
  assign PE_556_reset = reset;
  assign PE_556_io_data_2_sig_stat2trans = PENetwork_77_io_to_pes_6_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_556_io_data_1_in_valid = PENetwork_47_io_to_pes_6_in_valid; // @[pe.scala 264:34]
  assign PE_556_io_data_1_in_bits = PENetwork_47_io_to_pes_6_in_bits; // @[pe.scala 264:34]
  assign PE_556_io_data_0_in_valid = PENetwork_6_io_to_pes_25_in_valid; // @[pe.scala 264:34]
  assign PE_556_io_data_0_in_bits = PENetwork_6_io_to_pes_25_in_bits; // @[pe.scala 264:34]
  assign PE_557_clock = clock;
  assign PE_557_reset = reset;
  assign PE_557_io_data_2_sig_stat2trans = PENetwork_77_io_to_pes_7_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_557_io_data_1_in_valid = PENetwork_47_io_to_pes_7_in_valid; // @[pe.scala 264:34]
  assign PE_557_io_data_1_in_bits = PENetwork_47_io_to_pes_7_in_bits; // @[pe.scala 264:34]
  assign PE_557_io_data_0_in_valid = PENetwork_7_io_to_pes_25_in_valid; // @[pe.scala 264:34]
  assign PE_557_io_data_0_in_bits = PENetwork_7_io_to_pes_25_in_bits; // @[pe.scala 264:34]
  assign PE_558_clock = clock;
  assign PE_558_reset = reset;
  assign PE_558_io_data_2_sig_stat2trans = PENetwork_77_io_to_pes_8_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_558_io_data_1_in_valid = PENetwork_47_io_to_pes_8_in_valid; // @[pe.scala 264:34]
  assign PE_558_io_data_1_in_bits = PENetwork_47_io_to_pes_8_in_bits; // @[pe.scala 264:34]
  assign PE_558_io_data_0_in_valid = PENetwork_8_io_to_pes_25_in_valid; // @[pe.scala 264:34]
  assign PE_558_io_data_0_in_bits = PENetwork_8_io_to_pes_25_in_bits; // @[pe.scala 264:34]
  assign PE_559_clock = clock;
  assign PE_559_reset = reset;
  assign PE_559_io_data_2_sig_stat2trans = PENetwork_77_io_to_pes_9_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_559_io_data_1_in_valid = PENetwork_47_io_to_pes_9_in_valid; // @[pe.scala 264:34]
  assign PE_559_io_data_1_in_bits = PENetwork_47_io_to_pes_9_in_bits; // @[pe.scala 264:34]
  assign PE_559_io_data_0_in_valid = PENetwork_9_io_to_pes_25_in_valid; // @[pe.scala 264:34]
  assign PE_559_io_data_0_in_bits = PENetwork_9_io_to_pes_25_in_bits; // @[pe.scala 264:34]
  assign PE_560_clock = clock;
  assign PE_560_reset = reset;
  assign PE_560_io_data_2_sig_stat2trans = PENetwork_77_io_to_pes_10_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_560_io_data_1_in_valid = PENetwork_47_io_to_pes_10_in_valid; // @[pe.scala 264:34]
  assign PE_560_io_data_1_in_bits = PENetwork_47_io_to_pes_10_in_bits; // @[pe.scala 264:34]
  assign PE_560_io_data_0_in_valid = PENetwork_10_io_to_pes_25_in_valid; // @[pe.scala 264:34]
  assign PE_560_io_data_0_in_bits = PENetwork_10_io_to_pes_25_in_bits; // @[pe.scala 264:34]
  assign PE_561_clock = clock;
  assign PE_561_reset = reset;
  assign PE_561_io_data_2_sig_stat2trans = PENetwork_77_io_to_pes_11_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_561_io_data_1_in_valid = PENetwork_47_io_to_pes_11_in_valid; // @[pe.scala 264:34]
  assign PE_561_io_data_1_in_bits = PENetwork_47_io_to_pes_11_in_bits; // @[pe.scala 264:34]
  assign PE_561_io_data_0_in_valid = PENetwork_11_io_to_pes_25_in_valid; // @[pe.scala 264:34]
  assign PE_561_io_data_0_in_bits = PENetwork_11_io_to_pes_25_in_bits; // @[pe.scala 264:34]
  assign PE_562_clock = clock;
  assign PE_562_reset = reset;
  assign PE_562_io_data_2_sig_stat2trans = PENetwork_77_io_to_pes_12_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_562_io_data_1_in_valid = PENetwork_47_io_to_pes_12_in_valid; // @[pe.scala 264:34]
  assign PE_562_io_data_1_in_bits = PENetwork_47_io_to_pes_12_in_bits; // @[pe.scala 264:34]
  assign PE_562_io_data_0_in_valid = PENetwork_12_io_to_pes_25_in_valid; // @[pe.scala 264:34]
  assign PE_562_io_data_0_in_bits = PENetwork_12_io_to_pes_25_in_bits; // @[pe.scala 264:34]
  assign PE_563_clock = clock;
  assign PE_563_reset = reset;
  assign PE_563_io_data_2_sig_stat2trans = PENetwork_77_io_to_pes_13_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_563_io_data_1_in_valid = PENetwork_47_io_to_pes_13_in_valid; // @[pe.scala 264:34]
  assign PE_563_io_data_1_in_bits = PENetwork_47_io_to_pes_13_in_bits; // @[pe.scala 264:34]
  assign PE_563_io_data_0_in_valid = PENetwork_13_io_to_pes_25_in_valid; // @[pe.scala 264:34]
  assign PE_563_io_data_0_in_bits = PENetwork_13_io_to_pes_25_in_bits; // @[pe.scala 264:34]
  assign PE_564_clock = clock;
  assign PE_564_reset = reset;
  assign PE_564_io_data_2_sig_stat2trans = PENetwork_77_io_to_pes_14_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_564_io_data_1_in_valid = PENetwork_47_io_to_pes_14_in_valid; // @[pe.scala 264:34]
  assign PE_564_io_data_1_in_bits = PENetwork_47_io_to_pes_14_in_bits; // @[pe.scala 264:34]
  assign PE_564_io_data_0_in_valid = PENetwork_14_io_to_pes_25_in_valid; // @[pe.scala 264:34]
  assign PE_564_io_data_0_in_bits = PENetwork_14_io_to_pes_25_in_bits; // @[pe.scala 264:34]
  assign PE_565_clock = clock;
  assign PE_565_reset = reset;
  assign PE_565_io_data_2_sig_stat2trans = PENetwork_77_io_to_pes_15_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_565_io_data_1_in_valid = PENetwork_47_io_to_pes_15_in_valid; // @[pe.scala 264:34]
  assign PE_565_io_data_1_in_bits = PENetwork_47_io_to_pes_15_in_bits; // @[pe.scala 264:34]
  assign PE_565_io_data_0_in_valid = PENetwork_15_io_to_pes_25_in_valid; // @[pe.scala 264:34]
  assign PE_565_io_data_0_in_bits = PENetwork_15_io_to_pes_25_in_bits; // @[pe.scala 264:34]
  assign PE_566_clock = clock;
  assign PE_566_reset = reset;
  assign PE_566_io_data_2_sig_stat2trans = PENetwork_77_io_to_pes_16_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_566_io_data_1_in_valid = PENetwork_47_io_to_pes_16_in_valid; // @[pe.scala 264:34]
  assign PE_566_io_data_1_in_bits = PENetwork_47_io_to_pes_16_in_bits; // @[pe.scala 264:34]
  assign PE_566_io_data_0_in_valid = PENetwork_16_io_to_pes_25_in_valid; // @[pe.scala 264:34]
  assign PE_566_io_data_0_in_bits = PENetwork_16_io_to_pes_25_in_bits; // @[pe.scala 264:34]
  assign PE_567_clock = clock;
  assign PE_567_reset = reset;
  assign PE_567_io_data_2_sig_stat2trans = PENetwork_77_io_to_pes_17_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_567_io_data_1_in_valid = PENetwork_47_io_to_pes_17_in_valid; // @[pe.scala 264:34]
  assign PE_567_io_data_1_in_bits = PENetwork_47_io_to_pes_17_in_bits; // @[pe.scala 264:34]
  assign PE_567_io_data_0_in_valid = PENetwork_17_io_to_pes_25_in_valid; // @[pe.scala 264:34]
  assign PE_567_io_data_0_in_bits = PENetwork_17_io_to_pes_25_in_bits; // @[pe.scala 264:34]
  assign PE_568_clock = clock;
  assign PE_568_reset = reset;
  assign PE_568_io_data_2_sig_stat2trans = PENetwork_77_io_to_pes_18_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_568_io_data_1_in_valid = PENetwork_47_io_to_pes_18_in_valid; // @[pe.scala 264:34]
  assign PE_568_io_data_1_in_bits = PENetwork_47_io_to_pes_18_in_bits; // @[pe.scala 264:34]
  assign PE_568_io_data_0_in_valid = PENetwork_18_io_to_pes_25_in_valid; // @[pe.scala 264:34]
  assign PE_568_io_data_0_in_bits = PENetwork_18_io_to_pes_25_in_bits; // @[pe.scala 264:34]
  assign PE_569_clock = clock;
  assign PE_569_reset = reset;
  assign PE_569_io_data_2_sig_stat2trans = PENetwork_77_io_to_pes_19_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_569_io_data_1_in_valid = PENetwork_47_io_to_pes_19_in_valid; // @[pe.scala 264:34]
  assign PE_569_io_data_1_in_bits = PENetwork_47_io_to_pes_19_in_bits; // @[pe.scala 264:34]
  assign PE_569_io_data_0_in_valid = PENetwork_19_io_to_pes_25_in_valid; // @[pe.scala 264:34]
  assign PE_569_io_data_0_in_bits = PENetwork_19_io_to_pes_25_in_bits; // @[pe.scala 264:34]
  assign PE_570_clock = clock;
  assign PE_570_reset = reset;
  assign PE_570_io_data_2_sig_stat2trans = PENetwork_77_io_to_pes_20_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_570_io_data_1_in_valid = PENetwork_47_io_to_pes_20_in_valid; // @[pe.scala 264:34]
  assign PE_570_io_data_1_in_bits = PENetwork_47_io_to_pes_20_in_bits; // @[pe.scala 264:34]
  assign PE_570_io_data_0_in_valid = PENetwork_20_io_to_pes_25_in_valid; // @[pe.scala 264:34]
  assign PE_570_io_data_0_in_bits = PENetwork_20_io_to_pes_25_in_bits; // @[pe.scala 264:34]
  assign PE_571_clock = clock;
  assign PE_571_reset = reset;
  assign PE_571_io_data_2_sig_stat2trans = PENetwork_77_io_to_pes_21_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_571_io_data_1_in_valid = PENetwork_47_io_to_pes_21_in_valid; // @[pe.scala 264:34]
  assign PE_571_io_data_1_in_bits = PENetwork_47_io_to_pes_21_in_bits; // @[pe.scala 264:34]
  assign PE_571_io_data_0_in_valid = PENetwork_21_io_to_pes_25_in_valid; // @[pe.scala 264:34]
  assign PE_571_io_data_0_in_bits = PENetwork_21_io_to_pes_25_in_bits; // @[pe.scala 264:34]
  assign PE_572_clock = clock;
  assign PE_572_reset = reset;
  assign PE_572_io_data_2_sig_stat2trans = PENetwork_78_io_to_pes_0_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_572_io_data_1_in_valid = PENetwork_48_io_to_pes_0_in_valid; // @[pe.scala 264:34]
  assign PE_572_io_data_1_in_bits = PENetwork_48_io_to_pes_0_in_bits; // @[pe.scala 264:34]
  assign PE_572_io_data_0_in_valid = PENetwork_io_to_pes_26_in_valid; // @[pe.scala 264:34]
  assign PE_572_io_data_0_in_bits = PENetwork_io_to_pes_26_in_bits; // @[pe.scala 264:34]
  assign PE_573_clock = clock;
  assign PE_573_reset = reset;
  assign PE_573_io_data_2_sig_stat2trans = PENetwork_78_io_to_pes_1_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_573_io_data_1_in_valid = PENetwork_48_io_to_pes_1_in_valid; // @[pe.scala 264:34]
  assign PE_573_io_data_1_in_bits = PENetwork_48_io_to_pes_1_in_bits; // @[pe.scala 264:34]
  assign PE_573_io_data_0_in_valid = PENetwork_1_io_to_pes_26_in_valid; // @[pe.scala 264:34]
  assign PE_573_io_data_0_in_bits = PENetwork_1_io_to_pes_26_in_bits; // @[pe.scala 264:34]
  assign PE_574_clock = clock;
  assign PE_574_reset = reset;
  assign PE_574_io_data_2_sig_stat2trans = PENetwork_78_io_to_pes_2_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_574_io_data_1_in_valid = PENetwork_48_io_to_pes_2_in_valid; // @[pe.scala 264:34]
  assign PE_574_io_data_1_in_bits = PENetwork_48_io_to_pes_2_in_bits; // @[pe.scala 264:34]
  assign PE_574_io_data_0_in_valid = PENetwork_2_io_to_pes_26_in_valid; // @[pe.scala 264:34]
  assign PE_574_io_data_0_in_bits = PENetwork_2_io_to_pes_26_in_bits; // @[pe.scala 264:34]
  assign PE_575_clock = clock;
  assign PE_575_reset = reset;
  assign PE_575_io_data_2_sig_stat2trans = PENetwork_78_io_to_pes_3_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_575_io_data_1_in_valid = PENetwork_48_io_to_pes_3_in_valid; // @[pe.scala 264:34]
  assign PE_575_io_data_1_in_bits = PENetwork_48_io_to_pes_3_in_bits; // @[pe.scala 264:34]
  assign PE_575_io_data_0_in_valid = PENetwork_3_io_to_pes_26_in_valid; // @[pe.scala 264:34]
  assign PE_575_io_data_0_in_bits = PENetwork_3_io_to_pes_26_in_bits; // @[pe.scala 264:34]
  assign PE_576_clock = clock;
  assign PE_576_reset = reset;
  assign PE_576_io_data_2_sig_stat2trans = PENetwork_78_io_to_pes_4_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_576_io_data_1_in_valid = PENetwork_48_io_to_pes_4_in_valid; // @[pe.scala 264:34]
  assign PE_576_io_data_1_in_bits = PENetwork_48_io_to_pes_4_in_bits; // @[pe.scala 264:34]
  assign PE_576_io_data_0_in_valid = PENetwork_4_io_to_pes_26_in_valid; // @[pe.scala 264:34]
  assign PE_576_io_data_0_in_bits = PENetwork_4_io_to_pes_26_in_bits; // @[pe.scala 264:34]
  assign PE_577_clock = clock;
  assign PE_577_reset = reset;
  assign PE_577_io_data_2_sig_stat2trans = PENetwork_78_io_to_pes_5_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_577_io_data_1_in_valid = PENetwork_48_io_to_pes_5_in_valid; // @[pe.scala 264:34]
  assign PE_577_io_data_1_in_bits = PENetwork_48_io_to_pes_5_in_bits; // @[pe.scala 264:34]
  assign PE_577_io_data_0_in_valid = PENetwork_5_io_to_pes_26_in_valid; // @[pe.scala 264:34]
  assign PE_577_io_data_0_in_bits = PENetwork_5_io_to_pes_26_in_bits; // @[pe.scala 264:34]
  assign PE_578_clock = clock;
  assign PE_578_reset = reset;
  assign PE_578_io_data_2_sig_stat2trans = PENetwork_78_io_to_pes_6_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_578_io_data_1_in_valid = PENetwork_48_io_to_pes_6_in_valid; // @[pe.scala 264:34]
  assign PE_578_io_data_1_in_bits = PENetwork_48_io_to_pes_6_in_bits; // @[pe.scala 264:34]
  assign PE_578_io_data_0_in_valid = PENetwork_6_io_to_pes_26_in_valid; // @[pe.scala 264:34]
  assign PE_578_io_data_0_in_bits = PENetwork_6_io_to_pes_26_in_bits; // @[pe.scala 264:34]
  assign PE_579_clock = clock;
  assign PE_579_reset = reset;
  assign PE_579_io_data_2_sig_stat2trans = PENetwork_78_io_to_pes_7_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_579_io_data_1_in_valid = PENetwork_48_io_to_pes_7_in_valid; // @[pe.scala 264:34]
  assign PE_579_io_data_1_in_bits = PENetwork_48_io_to_pes_7_in_bits; // @[pe.scala 264:34]
  assign PE_579_io_data_0_in_valid = PENetwork_7_io_to_pes_26_in_valid; // @[pe.scala 264:34]
  assign PE_579_io_data_0_in_bits = PENetwork_7_io_to_pes_26_in_bits; // @[pe.scala 264:34]
  assign PE_580_clock = clock;
  assign PE_580_reset = reset;
  assign PE_580_io_data_2_sig_stat2trans = PENetwork_78_io_to_pes_8_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_580_io_data_1_in_valid = PENetwork_48_io_to_pes_8_in_valid; // @[pe.scala 264:34]
  assign PE_580_io_data_1_in_bits = PENetwork_48_io_to_pes_8_in_bits; // @[pe.scala 264:34]
  assign PE_580_io_data_0_in_valid = PENetwork_8_io_to_pes_26_in_valid; // @[pe.scala 264:34]
  assign PE_580_io_data_0_in_bits = PENetwork_8_io_to_pes_26_in_bits; // @[pe.scala 264:34]
  assign PE_581_clock = clock;
  assign PE_581_reset = reset;
  assign PE_581_io_data_2_sig_stat2trans = PENetwork_78_io_to_pes_9_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_581_io_data_1_in_valid = PENetwork_48_io_to_pes_9_in_valid; // @[pe.scala 264:34]
  assign PE_581_io_data_1_in_bits = PENetwork_48_io_to_pes_9_in_bits; // @[pe.scala 264:34]
  assign PE_581_io_data_0_in_valid = PENetwork_9_io_to_pes_26_in_valid; // @[pe.scala 264:34]
  assign PE_581_io_data_0_in_bits = PENetwork_9_io_to_pes_26_in_bits; // @[pe.scala 264:34]
  assign PE_582_clock = clock;
  assign PE_582_reset = reset;
  assign PE_582_io_data_2_sig_stat2trans = PENetwork_78_io_to_pes_10_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_582_io_data_1_in_valid = PENetwork_48_io_to_pes_10_in_valid; // @[pe.scala 264:34]
  assign PE_582_io_data_1_in_bits = PENetwork_48_io_to_pes_10_in_bits; // @[pe.scala 264:34]
  assign PE_582_io_data_0_in_valid = PENetwork_10_io_to_pes_26_in_valid; // @[pe.scala 264:34]
  assign PE_582_io_data_0_in_bits = PENetwork_10_io_to_pes_26_in_bits; // @[pe.scala 264:34]
  assign PE_583_clock = clock;
  assign PE_583_reset = reset;
  assign PE_583_io_data_2_sig_stat2trans = PENetwork_78_io_to_pes_11_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_583_io_data_1_in_valid = PENetwork_48_io_to_pes_11_in_valid; // @[pe.scala 264:34]
  assign PE_583_io_data_1_in_bits = PENetwork_48_io_to_pes_11_in_bits; // @[pe.scala 264:34]
  assign PE_583_io_data_0_in_valid = PENetwork_11_io_to_pes_26_in_valid; // @[pe.scala 264:34]
  assign PE_583_io_data_0_in_bits = PENetwork_11_io_to_pes_26_in_bits; // @[pe.scala 264:34]
  assign PE_584_clock = clock;
  assign PE_584_reset = reset;
  assign PE_584_io_data_2_sig_stat2trans = PENetwork_78_io_to_pes_12_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_584_io_data_1_in_valid = PENetwork_48_io_to_pes_12_in_valid; // @[pe.scala 264:34]
  assign PE_584_io_data_1_in_bits = PENetwork_48_io_to_pes_12_in_bits; // @[pe.scala 264:34]
  assign PE_584_io_data_0_in_valid = PENetwork_12_io_to_pes_26_in_valid; // @[pe.scala 264:34]
  assign PE_584_io_data_0_in_bits = PENetwork_12_io_to_pes_26_in_bits; // @[pe.scala 264:34]
  assign PE_585_clock = clock;
  assign PE_585_reset = reset;
  assign PE_585_io_data_2_sig_stat2trans = PENetwork_78_io_to_pes_13_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_585_io_data_1_in_valid = PENetwork_48_io_to_pes_13_in_valid; // @[pe.scala 264:34]
  assign PE_585_io_data_1_in_bits = PENetwork_48_io_to_pes_13_in_bits; // @[pe.scala 264:34]
  assign PE_585_io_data_0_in_valid = PENetwork_13_io_to_pes_26_in_valid; // @[pe.scala 264:34]
  assign PE_585_io_data_0_in_bits = PENetwork_13_io_to_pes_26_in_bits; // @[pe.scala 264:34]
  assign PE_586_clock = clock;
  assign PE_586_reset = reset;
  assign PE_586_io_data_2_sig_stat2trans = PENetwork_78_io_to_pes_14_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_586_io_data_1_in_valid = PENetwork_48_io_to_pes_14_in_valid; // @[pe.scala 264:34]
  assign PE_586_io_data_1_in_bits = PENetwork_48_io_to_pes_14_in_bits; // @[pe.scala 264:34]
  assign PE_586_io_data_0_in_valid = PENetwork_14_io_to_pes_26_in_valid; // @[pe.scala 264:34]
  assign PE_586_io_data_0_in_bits = PENetwork_14_io_to_pes_26_in_bits; // @[pe.scala 264:34]
  assign PE_587_clock = clock;
  assign PE_587_reset = reset;
  assign PE_587_io_data_2_sig_stat2trans = PENetwork_78_io_to_pes_15_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_587_io_data_1_in_valid = PENetwork_48_io_to_pes_15_in_valid; // @[pe.scala 264:34]
  assign PE_587_io_data_1_in_bits = PENetwork_48_io_to_pes_15_in_bits; // @[pe.scala 264:34]
  assign PE_587_io_data_0_in_valid = PENetwork_15_io_to_pes_26_in_valid; // @[pe.scala 264:34]
  assign PE_587_io_data_0_in_bits = PENetwork_15_io_to_pes_26_in_bits; // @[pe.scala 264:34]
  assign PE_588_clock = clock;
  assign PE_588_reset = reset;
  assign PE_588_io_data_2_sig_stat2trans = PENetwork_78_io_to_pes_16_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_588_io_data_1_in_valid = PENetwork_48_io_to_pes_16_in_valid; // @[pe.scala 264:34]
  assign PE_588_io_data_1_in_bits = PENetwork_48_io_to_pes_16_in_bits; // @[pe.scala 264:34]
  assign PE_588_io_data_0_in_valid = PENetwork_16_io_to_pes_26_in_valid; // @[pe.scala 264:34]
  assign PE_588_io_data_0_in_bits = PENetwork_16_io_to_pes_26_in_bits; // @[pe.scala 264:34]
  assign PE_589_clock = clock;
  assign PE_589_reset = reset;
  assign PE_589_io_data_2_sig_stat2trans = PENetwork_78_io_to_pes_17_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_589_io_data_1_in_valid = PENetwork_48_io_to_pes_17_in_valid; // @[pe.scala 264:34]
  assign PE_589_io_data_1_in_bits = PENetwork_48_io_to_pes_17_in_bits; // @[pe.scala 264:34]
  assign PE_589_io_data_0_in_valid = PENetwork_17_io_to_pes_26_in_valid; // @[pe.scala 264:34]
  assign PE_589_io_data_0_in_bits = PENetwork_17_io_to_pes_26_in_bits; // @[pe.scala 264:34]
  assign PE_590_clock = clock;
  assign PE_590_reset = reset;
  assign PE_590_io_data_2_sig_stat2trans = PENetwork_78_io_to_pes_18_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_590_io_data_1_in_valid = PENetwork_48_io_to_pes_18_in_valid; // @[pe.scala 264:34]
  assign PE_590_io_data_1_in_bits = PENetwork_48_io_to_pes_18_in_bits; // @[pe.scala 264:34]
  assign PE_590_io_data_0_in_valid = PENetwork_18_io_to_pes_26_in_valid; // @[pe.scala 264:34]
  assign PE_590_io_data_0_in_bits = PENetwork_18_io_to_pes_26_in_bits; // @[pe.scala 264:34]
  assign PE_591_clock = clock;
  assign PE_591_reset = reset;
  assign PE_591_io_data_2_sig_stat2trans = PENetwork_78_io_to_pes_19_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_591_io_data_1_in_valid = PENetwork_48_io_to_pes_19_in_valid; // @[pe.scala 264:34]
  assign PE_591_io_data_1_in_bits = PENetwork_48_io_to_pes_19_in_bits; // @[pe.scala 264:34]
  assign PE_591_io_data_0_in_valid = PENetwork_19_io_to_pes_26_in_valid; // @[pe.scala 264:34]
  assign PE_591_io_data_0_in_bits = PENetwork_19_io_to_pes_26_in_bits; // @[pe.scala 264:34]
  assign PE_592_clock = clock;
  assign PE_592_reset = reset;
  assign PE_592_io_data_2_sig_stat2trans = PENetwork_78_io_to_pes_20_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_592_io_data_1_in_valid = PENetwork_48_io_to_pes_20_in_valid; // @[pe.scala 264:34]
  assign PE_592_io_data_1_in_bits = PENetwork_48_io_to_pes_20_in_bits; // @[pe.scala 264:34]
  assign PE_592_io_data_0_in_valid = PENetwork_20_io_to_pes_26_in_valid; // @[pe.scala 264:34]
  assign PE_592_io_data_0_in_bits = PENetwork_20_io_to_pes_26_in_bits; // @[pe.scala 264:34]
  assign PE_593_clock = clock;
  assign PE_593_reset = reset;
  assign PE_593_io_data_2_sig_stat2trans = PENetwork_78_io_to_pes_21_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_593_io_data_1_in_valid = PENetwork_48_io_to_pes_21_in_valid; // @[pe.scala 264:34]
  assign PE_593_io_data_1_in_bits = PENetwork_48_io_to_pes_21_in_bits; // @[pe.scala 264:34]
  assign PE_593_io_data_0_in_valid = PENetwork_21_io_to_pes_26_in_valid; // @[pe.scala 264:34]
  assign PE_593_io_data_0_in_bits = PENetwork_21_io_to_pes_26_in_bits; // @[pe.scala 264:34]
  assign PE_594_clock = clock;
  assign PE_594_reset = reset;
  assign PE_594_io_data_2_sig_stat2trans = PENetwork_79_io_to_pes_0_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_594_io_data_1_in_valid = PENetwork_49_io_to_pes_0_in_valid; // @[pe.scala 264:34]
  assign PE_594_io_data_1_in_bits = PENetwork_49_io_to_pes_0_in_bits; // @[pe.scala 264:34]
  assign PE_594_io_data_0_in_valid = PENetwork_io_to_pes_27_in_valid; // @[pe.scala 264:34]
  assign PE_594_io_data_0_in_bits = PENetwork_io_to_pes_27_in_bits; // @[pe.scala 264:34]
  assign PE_595_clock = clock;
  assign PE_595_reset = reset;
  assign PE_595_io_data_2_sig_stat2trans = PENetwork_79_io_to_pes_1_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_595_io_data_1_in_valid = PENetwork_49_io_to_pes_1_in_valid; // @[pe.scala 264:34]
  assign PE_595_io_data_1_in_bits = PENetwork_49_io_to_pes_1_in_bits; // @[pe.scala 264:34]
  assign PE_595_io_data_0_in_valid = PENetwork_1_io_to_pes_27_in_valid; // @[pe.scala 264:34]
  assign PE_595_io_data_0_in_bits = PENetwork_1_io_to_pes_27_in_bits; // @[pe.scala 264:34]
  assign PE_596_clock = clock;
  assign PE_596_reset = reset;
  assign PE_596_io_data_2_sig_stat2trans = PENetwork_79_io_to_pes_2_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_596_io_data_1_in_valid = PENetwork_49_io_to_pes_2_in_valid; // @[pe.scala 264:34]
  assign PE_596_io_data_1_in_bits = PENetwork_49_io_to_pes_2_in_bits; // @[pe.scala 264:34]
  assign PE_596_io_data_0_in_valid = PENetwork_2_io_to_pes_27_in_valid; // @[pe.scala 264:34]
  assign PE_596_io_data_0_in_bits = PENetwork_2_io_to_pes_27_in_bits; // @[pe.scala 264:34]
  assign PE_597_clock = clock;
  assign PE_597_reset = reset;
  assign PE_597_io_data_2_sig_stat2trans = PENetwork_79_io_to_pes_3_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_597_io_data_1_in_valid = PENetwork_49_io_to_pes_3_in_valid; // @[pe.scala 264:34]
  assign PE_597_io_data_1_in_bits = PENetwork_49_io_to_pes_3_in_bits; // @[pe.scala 264:34]
  assign PE_597_io_data_0_in_valid = PENetwork_3_io_to_pes_27_in_valid; // @[pe.scala 264:34]
  assign PE_597_io_data_0_in_bits = PENetwork_3_io_to_pes_27_in_bits; // @[pe.scala 264:34]
  assign PE_598_clock = clock;
  assign PE_598_reset = reset;
  assign PE_598_io_data_2_sig_stat2trans = PENetwork_79_io_to_pes_4_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_598_io_data_1_in_valid = PENetwork_49_io_to_pes_4_in_valid; // @[pe.scala 264:34]
  assign PE_598_io_data_1_in_bits = PENetwork_49_io_to_pes_4_in_bits; // @[pe.scala 264:34]
  assign PE_598_io_data_0_in_valid = PENetwork_4_io_to_pes_27_in_valid; // @[pe.scala 264:34]
  assign PE_598_io_data_0_in_bits = PENetwork_4_io_to_pes_27_in_bits; // @[pe.scala 264:34]
  assign PE_599_clock = clock;
  assign PE_599_reset = reset;
  assign PE_599_io_data_2_sig_stat2trans = PENetwork_79_io_to_pes_5_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_599_io_data_1_in_valid = PENetwork_49_io_to_pes_5_in_valid; // @[pe.scala 264:34]
  assign PE_599_io_data_1_in_bits = PENetwork_49_io_to_pes_5_in_bits; // @[pe.scala 264:34]
  assign PE_599_io_data_0_in_valid = PENetwork_5_io_to_pes_27_in_valid; // @[pe.scala 264:34]
  assign PE_599_io_data_0_in_bits = PENetwork_5_io_to_pes_27_in_bits; // @[pe.scala 264:34]
  assign PE_600_clock = clock;
  assign PE_600_reset = reset;
  assign PE_600_io_data_2_sig_stat2trans = PENetwork_79_io_to_pes_6_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_600_io_data_1_in_valid = PENetwork_49_io_to_pes_6_in_valid; // @[pe.scala 264:34]
  assign PE_600_io_data_1_in_bits = PENetwork_49_io_to_pes_6_in_bits; // @[pe.scala 264:34]
  assign PE_600_io_data_0_in_valid = PENetwork_6_io_to_pes_27_in_valid; // @[pe.scala 264:34]
  assign PE_600_io_data_0_in_bits = PENetwork_6_io_to_pes_27_in_bits; // @[pe.scala 264:34]
  assign PE_601_clock = clock;
  assign PE_601_reset = reset;
  assign PE_601_io_data_2_sig_stat2trans = PENetwork_79_io_to_pes_7_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_601_io_data_1_in_valid = PENetwork_49_io_to_pes_7_in_valid; // @[pe.scala 264:34]
  assign PE_601_io_data_1_in_bits = PENetwork_49_io_to_pes_7_in_bits; // @[pe.scala 264:34]
  assign PE_601_io_data_0_in_valid = PENetwork_7_io_to_pes_27_in_valid; // @[pe.scala 264:34]
  assign PE_601_io_data_0_in_bits = PENetwork_7_io_to_pes_27_in_bits; // @[pe.scala 264:34]
  assign PE_602_clock = clock;
  assign PE_602_reset = reset;
  assign PE_602_io_data_2_sig_stat2trans = PENetwork_79_io_to_pes_8_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_602_io_data_1_in_valid = PENetwork_49_io_to_pes_8_in_valid; // @[pe.scala 264:34]
  assign PE_602_io_data_1_in_bits = PENetwork_49_io_to_pes_8_in_bits; // @[pe.scala 264:34]
  assign PE_602_io_data_0_in_valid = PENetwork_8_io_to_pes_27_in_valid; // @[pe.scala 264:34]
  assign PE_602_io_data_0_in_bits = PENetwork_8_io_to_pes_27_in_bits; // @[pe.scala 264:34]
  assign PE_603_clock = clock;
  assign PE_603_reset = reset;
  assign PE_603_io_data_2_sig_stat2trans = PENetwork_79_io_to_pes_9_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_603_io_data_1_in_valid = PENetwork_49_io_to_pes_9_in_valid; // @[pe.scala 264:34]
  assign PE_603_io_data_1_in_bits = PENetwork_49_io_to_pes_9_in_bits; // @[pe.scala 264:34]
  assign PE_603_io_data_0_in_valid = PENetwork_9_io_to_pes_27_in_valid; // @[pe.scala 264:34]
  assign PE_603_io_data_0_in_bits = PENetwork_9_io_to_pes_27_in_bits; // @[pe.scala 264:34]
  assign PE_604_clock = clock;
  assign PE_604_reset = reset;
  assign PE_604_io_data_2_sig_stat2trans = PENetwork_79_io_to_pes_10_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_604_io_data_1_in_valid = PENetwork_49_io_to_pes_10_in_valid; // @[pe.scala 264:34]
  assign PE_604_io_data_1_in_bits = PENetwork_49_io_to_pes_10_in_bits; // @[pe.scala 264:34]
  assign PE_604_io_data_0_in_valid = PENetwork_10_io_to_pes_27_in_valid; // @[pe.scala 264:34]
  assign PE_604_io_data_0_in_bits = PENetwork_10_io_to_pes_27_in_bits; // @[pe.scala 264:34]
  assign PE_605_clock = clock;
  assign PE_605_reset = reset;
  assign PE_605_io_data_2_sig_stat2trans = PENetwork_79_io_to_pes_11_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_605_io_data_1_in_valid = PENetwork_49_io_to_pes_11_in_valid; // @[pe.scala 264:34]
  assign PE_605_io_data_1_in_bits = PENetwork_49_io_to_pes_11_in_bits; // @[pe.scala 264:34]
  assign PE_605_io_data_0_in_valid = PENetwork_11_io_to_pes_27_in_valid; // @[pe.scala 264:34]
  assign PE_605_io_data_0_in_bits = PENetwork_11_io_to_pes_27_in_bits; // @[pe.scala 264:34]
  assign PE_606_clock = clock;
  assign PE_606_reset = reset;
  assign PE_606_io_data_2_sig_stat2trans = PENetwork_79_io_to_pes_12_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_606_io_data_1_in_valid = PENetwork_49_io_to_pes_12_in_valid; // @[pe.scala 264:34]
  assign PE_606_io_data_1_in_bits = PENetwork_49_io_to_pes_12_in_bits; // @[pe.scala 264:34]
  assign PE_606_io_data_0_in_valid = PENetwork_12_io_to_pes_27_in_valid; // @[pe.scala 264:34]
  assign PE_606_io_data_0_in_bits = PENetwork_12_io_to_pes_27_in_bits; // @[pe.scala 264:34]
  assign PE_607_clock = clock;
  assign PE_607_reset = reset;
  assign PE_607_io_data_2_sig_stat2trans = PENetwork_79_io_to_pes_13_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_607_io_data_1_in_valid = PENetwork_49_io_to_pes_13_in_valid; // @[pe.scala 264:34]
  assign PE_607_io_data_1_in_bits = PENetwork_49_io_to_pes_13_in_bits; // @[pe.scala 264:34]
  assign PE_607_io_data_0_in_valid = PENetwork_13_io_to_pes_27_in_valid; // @[pe.scala 264:34]
  assign PE_607_io_data_0_in_bits = PENetwork_13_io_to_pes_27_in_bits; // @[pe.scala 264:34]
  assign PE_608_clock = clock;
  assign PE_608_reset = reset;
  assign PE_608_io_data_2_sig_stat2trans = PENetwork_79_io_to_pes_14_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_608_io_data_1_in_valid = PENetwork_49_io_to_pes_14_in_valid; // @[pe.scala 264:34]
  assign PE_608_io_data_1_in_bits = PENetwork_49_io_to_pes_14_in_bits; // @[pe.scala 264:34]
  assign PE_608_io_data_0_in_valid = PENetwork_14_io_to_pes_27_in_valid; // @[pe.scala 264:34]
  assign PE_608_io_data_0_in_bits = PENetwork_14_io_to_pes_27_in_bits; // @[pe.scala 264:34]
  assign PE_609_clock = clock;
  assign PE_609_reset = reset;
  assign PE_609_io_data_2_sig_stat2trans = PENetwork_79_io_to_pes_15_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_609_io_data_1_in_valid = PENetwork_49_io_to_pes_15_in_valid; // @[pe.scala 264:34]
  assign PE_609_io_data_1_in_bits = PENetwork_49_io_to_pes_15_in_bits; // @[pe.scala 264:34]
  assign PE_609_io_data_0_in_valid = PENetwork_15_io_to_pes_27_in_valid; // @[pe.scala 264:34]
  assign PE_609_io_data_0_in_bits = PENetwork_15_io_to_pes_27_in_bits; // @[pe.scala 264:34]
  assign PE_610_clock = clock;
  assign PE_610_reset = reset;
  assign PE_610_io_data_2_sig_stat2trans = PENetwork_79_io_to_pes_16_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_610_io_data_1_in_valid = PENetwork_49_io_to_pes_16_in_valid; // @[pe.scala 264:34]
  assign PE_610_io_data_1_in_bits = PENetwork_49_io_to_pes_16_in_bits; // @[pe.scala 264:34]
  assign PE_610_io_data_0_in_valid = PENetwork_16_io_to_pes_27_in_valid; // @[pe.scala 264:34]
  assign PE_610_io_data_0_in_bits = PENetwork_16_io_to_pes_27_in_bits; // @[pe.scala 264:34]
  assign PE_611_clock = clock;
  assign PE_611_reset = reset;
  assign PE_611_io_data_2_sig_stat2trans = PENetwork_79_io_to_pes_17_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_611_io_data_1_in_valid = PENetwork_49_io_to_pes_17_in_valid; // @[pe.scala 264:34]
  assign PE_611_io_data_1_in_bits = PENetwork_49_io_to_pes_17_in_bits; // @[pe.scala 264:34]
  assign PE_611_io_data_0_in_valid = PENetwork_17_io_to_pes_27_in_valid; // @[pe.scala 264:34]
  assign PE_611_io_data_0_in_bits = PENetwork_17_io_to_pes_27_in_bits; // @[pe.scala 264:34]
  assign PE_612_clock = clock;
  assign PE_612_reset = reset;
  assign PE_612_io_data_2_sig_stat2trans = PENetwork_79_io_to_pes_18_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_612_io_data_1_in_valid = PENetwork_49_io_to_pes_18_in_valid; // @[pe.scala 264:34]
  assign PE_612_io_data_1_in_bits = PENetwork_49_io_to_pes_18_in_bits; // @[pe.scala 264:34]
  assign PE_612_io_data_0_in_valid = PENetwork_18_io_to_pes_27_in_valid; // @[pe.scala 264:34]
  assign PE_612_io_data_0_in_bits = PENetwork_18_io_to_pes_27_in_bits; // @[pe.scala 264:34]
  assign PE_613_clock = clock;
  assign PE_613_reset = reset;
  assign PE_613_io_data_2_sig_stat2trans = PENetwork_79_io_to_pes_19_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_613_io_data_1_in_valid = PENetwork_49_io_to_pes_19_in_valid; // @[pe.scala 264:34]
  assign PE_613_io_data_1_in_bits = PENetwork_49_io_to_pes_19_in_bits; // @[pe.scala 264:34]
  assign PE_613_io_data_0_in_valid = PENetwork_19_io_to_pes_27_in_valid; // @[pe.scala 264:34]
  assign PE_613_io_data_0_in_bits = PENetwork_19_io_to_pes_27_in_bits; // @[pe.scala 264:34]
  assign PE_614_clock = clock;
  assign PE_614_reset = reset;
  assign PE_614_io_data_2_sig_stat2trans = PENetwork_79_io_to_pes_20_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_614_io_data_1_in_valid = PENetwork_49_io_to_pes_20_in_valid; // @[pe.scala 264:34]
  assign PE_614_io_data_1_in_bits = PENetwork_49_io_to_pes_20_in_bits; // @[pe.scala 264:34]
  assign PE_614_io_data_0_in_valid = PENetwork_20_io_to_pes_27_in_valid; // @[pe.scala 264:34]
  assign PE_614_io_data_0_in_bits = PENetwork_20_io_to_pes_27_in_bits; // @[pe.scala 264:34]
  assign PE_615_clock = clock;
  assign PE_615_reset = reset;
  assign PE_615_io_data_2_sig_stat2trans = PENetwork_79_io_to_pes_21_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_615_io_data_1_in_valid = PENetwork_49_io_to_pes_21_in_valid; // @[pe.scala 264:34]
  assign PE_615_io_data_1_in_bits = PENetwork_49_io_to_pes_21_in_bits; // @[pe.scala 264:34]
  assign PE_615_io_data_0_in_valid = PENetwork_21_io_to_pes_27_in_valid; // @[pe.scala 264:34]
  assign PE_615_io_data_0_in_bits = PENetwork_21_io_to_pes_27_in_bits; // @[pe.scala 264:34]
  assign PE_616_clock = clock;
  assign PE_616_reset = reset;
  assign PE_616_io_data_2_sig_stat2trans = PENetwork_80_io_to_pes_0_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_616_io_data_1_in_valid = PENetwork_50_io_to_pes_0_in_valid; // @[pe.scala 264:34]
  assign PE_616_io_data_1_in_bits = PENetwork_50_io_to_pes_0_in_bits; // @[pe.scala 264:34]
  assign PE_616_io_data_0_in_valid = PENetwork_io_to_pes_28_in_valid; // @[pe.scala 264:34]
  assign PE_616_io_data_0_in_bits = PENetwork_io_to_pes_28_in_bits; // @[pe.scala 264:34]
  assign PE_617_clock = clock;
  assign PE_617_reset = reset;
  assign PE_617_io_data_2_sig_stat2trans = PENetwork_80_io_to_pes_1_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_617_io_data_1_in_valid = PENetwork_50_io_to_pes_1_in_valid; // @[pe.scala 264:34]
  assign PE_617_io_data_1_in_bits = PENetwork_50_io_to_pes_1_in_bits; // @[pe.scala 264:34]
  assign PE_617_io_data_0_in_valid = PENetwork_1_io_to_pes_28_in_valid; // @[pe.scala 264:34]
  assign PE_617_io_data_0_in_bits = PENetwork_1_io_to_pes_28_in_bits; // @[pe.scala 264:34]
  assign PE_618_clock = clock;
  assign PE_618_reset = reset;
  assign PE_618_io_data_2_sig_stat2trans = PENetwork_80_io_to_pes_2_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_618_io_data_1_in_valid = PENetwork_50_io_to_pes_2_in_valid; // @[pe.scala 264:34]
  assign PE_618_io_data_1_in_bits = PENetwork_50_io_to_pes_2_in_bits; // @[pe.scala 264:34]
  assign PE_618_io_data_0_in_valid = PENetwork_2_io_to_pes_28_in_valid; // @[pe.scala 264:34]
  assign PE_618_io_data_0_in_bits = PENetwork_2_io_to_pes_28_in_bits; // @[pe.scala 264:34]
  assign PE_619_clock = clock;
  assign PE_619_reset = reset;
  assign PE_619_io_data_2_sig_stat2trans = PENetwork_80_io_to_pes_3_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_619_io_data_1_in_valid = PENetwork_50_io_to_pes_3_in_valid; // @[pe.scala 264:34]
  assign PE_619_io_data_1_in_bits = PENetwork_50_io_to_pes_3_in_bits; // @[pe.scala 264:34]
  assign PE_619_io_data_0_in_valid = PENetwork_3_io_to_pes_28_in_valid; // @[pe.scala 264:34]
  assign PE_619_io_data_0_in_bits = PENetwork_3_io_to_pes_28_in_bits; // @[pe.scala 264:34]
  assign PE_620_clock = clock;
  assign PE_620_reset = reset;
  assign PE_620_io_data_2_sig_stat2trans = PENetwork_80_io_to_pes_4_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_620_io_data_1_in_valid = PENetwork_50_io_to_pes_4_in_valid; // @[pe.scala 264:34]
  assign PE_620_io_data_1_in_bits = PENetwork_50_io_to_pes_4_in_bits; // @[pe.scala 264:34]
  assign PE_620_io_data_0_in_valid = PENetwork_4_io_to_pes_28_in_valid; // @[pe.scala 264:34]
  assign PE_620_io_data_0_in_bits = PENetwork_4_io_to_pes_28_in_bits; // @[pe.scala 264:34]
  assign PE_621_clock = clock;
  assign PE_621_reset = reset;
  assign PE_621_io_data_2_sig_stat2trans = PENetwork_80_io_to_pes_5_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_621_io_data_1_in_valid = PENetwork_50_io_to_pes_5_in_valid; // @[pe.scala 264:34]
  assign PE_621_io_data_1_in_bits = PENetwork_50_io_to_pes_5_in_bits; // @[pe.scala 264:34]
  assign PE_621_io_data_0_in_valid = PENetwork_5_io_to_pes_28_in_valid; // @[pe.scala 264:34]
  assign PE_621_io_data_0_in_bits = PENetwork_5_io_to_pes_28_in_bits; // @[pe.scala 264:34]
  assign PE_622_clock = clock;
  assign PE_622_reset = reset;
  assign PE_622_io_data_2_sig_stat2trans = PENetwork_80_io_to_pes_6_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_622_io_data_1_in_valid = PENetwork_50_io_to_pes_6_in_valid; // @[pe.scala 264:34]
  assign PE_622_io_data_1_in_bits = PENetwork_50_io_to_pes_6_in_bits; // @[pe.scala 264:34]
  assign PE_622_io_data_0_in_valid = PENetwork_6_io_to_pes_28_in_valid; // @[pe.scala 264:34]
  assign PE_622_io_data_0_in_bits = PENetwork_6_io_to_pes_28_in_bits; // @[pe.scala 264:34]
  assign PE_623_clock = clock;
  assign PE_623_reset = reset;
  assign PE_623_io_data_2_sig_stat2trans = PENetwork_80_io_to_pes_7_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_623_io_data_1_in_valid = PENetwork_50_io_to_pes_7_in_valid; // @[pe.scala 264:34]
  assign PE_623_io_data_1_in_bits = PENetwork_50_io_to_pes_7_in_bits; // @[pe.scala 264:34]
  assign PE_623_io_data_0_in_valid = PENetwork_7_io_to_pes_28_in_valid; // @[pe.scala 264:34]
  assign PE_623_io_data_0_in_bits = PENetwork_7_io_to_pes_28_in_bits; // @[pe.scala 264:34]
  assign PE_624_clock = clock;
  assign PE_624_reset = reset;
  assign PE_624_io_data_2_sig_stat2trans = PENetwork_80_io_to_pes_8_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_624_io_data_1_in_valid = PENetwork_50_io_to_pes_8_in_valid; // @[pe.scala 264:34]
  assign PE_624_io_data_1_in_bits = PENetwork_50_io_to_pes_8_in_bits; // @[pe.scala 264:34]
  assign PE_624_io_data_0_in_valid = PENetwork_8_io_to_pes_28_in_valid; // @[pe.scala 264:34]
  assign PE_624_io_data_0_in_bits = PENetwork_8_io_to_pes_28_in_bits; // @[pe.scala 264:34]
  assign PE_625_clock = clock;
  assign PE_625_reset = reset;
  assign PE_625_io_data_2_sig_stat2trans = PENetwork_80_io_to_pes_9_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_625_io_data_1_in_valid = PENetwork_50_io_to_pes_9_in_valid; // @[pe.scala 264:34]
  assign PE_625_io_data_1_in_bits = PENetwork_50_io_to_pes_9_in_bits; // @[pe.scala 264:34]
  assign PE_625_io_data_0_in_valid = PENetwork_9_io_to_pes_28_in_valid; // @[pe.scala 264:34]
  assign PE_625_io_data_0_in_bits = PENetwork_9_io_to_pes_28_in_bits; // @[pe.scala 264:34]
  assign PE_626_clock = clock;
  assign PE_626_reset = reset;
  assign PE_626_io_data_2_sig_stat2trans = PENetwork_80_io_to_pes_10_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_626_io_data_1_in_valid = PENetwork_50_io_to_pes_10_in_valid; // @[pe.scala 264:34]
  assign PE_626_io_data_1_in_bits = PENetwork_50_io_to_pes_10_in_bits; // @[pe.scala 264:34]
  assign PE_626_io_data_0_in_valid = PENetwork_10_io_to_pes_28_in_valid; // @[pe.scala 264:34]
  assign PE_626_io_data_0_in_bits = PENetwork_10_io_to_pes_28_in_bits; // @[pe.scala 264:34]
  assign PE_627_clock = clock;
  assign PE_627_reset = reset;
  assign PE_627_io_data_2_sig_stat2trans = PENetwork_80_io_to_pes_11_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_627_io_data_1_in_valid = PENetwork_50_io_to_pes_11_in_valid; // @[pe.scala 264:34]
  assign PE_627_io_data_1_in_bits = PENetwork_50_io_to_pes_11_in_bits; // @[pe.scala 264:34]
  assign PE_627_io_data_0_in_valid = PENetwork_11_io_to_pes_28_in_valid; // @[pe.scala 264:34]
  assign PE_627_io_data_0_in_bits = PENetwork_11_io_to_pes_28_in_bits; // @[pe.scala 264:34]
  assign PE_628_clock = clock;
  assign PE_628_reset = reset;
  assign PE_628_io_data_2_sig_stat2trans = PENetwork_80_io_to_pes_12_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_628_io_data_1_in_valid = PENetwork_50_io_to_pes_12_in_valid; // @[pe.scala 264:34]
  assign PE_628_io_data_1_in_bits = PENetwork_50_io_to_pes_12_in_bits; // @[pe.scala 264:34]
  assign PE_628_io_data_0_in_valid = PENetwork_12_io_to_pes_28_in_valid; // @[pe.scala 264:34]
  assign PE_628_io_data_0_in_bits = PENetwork_12_io_to_pes_28_in_bits; // @[pe.scala 264:34]
  assign PE_629_clock = clock;
  assign PE_629_reset = reset;
  assign PE_629_io_data_2_sig_stat2trans = PENetwork_80_io_to_pes_13_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_629_io_data_1_in_valid = PENetwork_50_io_to_pes_13_in_valid; // @[pe.scala 264:34]
  assign PE_629_io_data_1_in_bits = PENetwork_50_io_to_pes_13_in_bits; // @[pe.scala 264:34]
  assign PE_629_io_data_0_in_valid = PENetwork_13_io_to_pes_28_in_valid; // @[pe.scala 264:34]
  assign PE_629_io_data_0_in_bits = PENetwork_13_io_to_pes_28_in_bits; // @[pe.scala 264:34]
  assign PE_630_clock = clock;
  assign PE_630_reset = reset;
  assign PE_630_io_data_2_sig_stat2trans = PENetwork_80_io_to_pes_14_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_630_io_data_1_in_valid = PENetwork_50_io_to_pes_14_in_valid; // @[pe.scala 264:34]
  assign PE_630_io_data_1_in_bits = PENetwork_50_io_to_pes_14_in_bits; // @[pe.scala 264:34]
  assign PE_630_io_data_0_in_valid = PENetwork_14_io_to_pes_28_in_valid; // @[pe.scala 264:34]
  assign PE_630_io_data_0_in_bits = PENetwork_14_io_to_pes_28_in_bits; // @[pe.scala 264:34]
  assign PE_631_clock = clock;
  assign PE_631_reset = reset;
  assign PE_631_io_data_2_sig_stat2trans = PENetwork_80_io_to_pes_15_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_631_io_data_1_in_valid = PENetwork_50_io_to_pes_15_in_valid; // @[pe.scala 264:34]
  assign PE_631_io_data_1_in_bits = PENetwork_50_io_to_pes_15_in_bits; // @[pe.scala 264:34]
  assign PE_631_io_data_0_in_valid = PENetwork_15_io_to_pes_28_in_valid; // @[pe.scala 264:34]
  assign PE_631_io_data_0_in_bits = PENetwork_15_io_to_pes_28_in_bits; // @[pe.scala 264:34]
  assign PE_632_clock = clock;
  assign PE_632_reset = reset;
  assign PE_632_io_data_2_sig_stat2trans = PENetwork_80_io_to_pes_16_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_632_io_data_1_in_valid = PENetwork_50_io_to_pes_16_in_valid; // @[pe.scala 264:34]
  assign PE_632_io_data_1_in_bits = PENetwork_50_io_to_pes_16_in_bits; // @[pe.scala 264:34]
  assign PE_632_io_data_0_in_valid = PENetwork_16_io_to_pes_28_in_valid; // @[pe.scala 264:34]
  assign PE_632_io_data_0_in_bits = PENetwork_16_io_to_pes_28_in_bits; // @[pe.scala 264:34]
  assign PE_633_clock = clock;
  assign PE_633_reset = reset;
  assign PE_633_io_data_2_sig_stat2trans = PENetwork_80_io_to_pes_17_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_633_io_data_1_in_valid = PENetwork_50_io_to_pes_17_in_valid; // @[pe.scala 264:34]
  assign PE_633_io_data_1_in_bits = PENetwork_50_io_to_pes_17_in_bits; // @[pe.scala 264:34]
  assign PE_633_io_data_0_in_valid = PENetwork_17_io_to_pes_28_in_valid; // @[pe.scala 264:34]
  assign PE_633_io_data_0_in_bits = PENetwork_17_io_to_pes_28_in_bits; // @[pe.scala 264:34]
  assign PE_634_clock = clock;
  assign PE_634_reset = reset;
  assign PE_634_io_data_2_sig_stat2trans = PENetwork_80_io_to_pes_18_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_634_io_data_1_in_valid = PENetwork_50_io_to_pes_18_in_valid; // @[pe.scala 264:34]
  assign PE_634_io_data_1_in_bits = PENetwork_50_io_to_pes_18_in_bits; // @[pe.scala 264:34]
  assign PE_634_io_data_0_in_valid = PENetwork_18_io_to_pes_28_in_valid; // @[pe.scala 264:34]
  assign PE_634_io_data_0_in_bits = PENetwork_18_io_to_pes_28_in_bits; // @[pe.scala 264:34]
  assign PE_635_clock = clock;
  assign PE_635_reset = reset;
  assign PE_635_io_data_2_sig_stat2trans = PENetwork_80_io_to_pes_19_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_635_io_data_1_in_valid = PENetwork_50_io_to_pes_19_in_valid; // @[pe.scala 264:34]
  assign PE_635_io_data_1_in_bits = PENetwork_50_io_to_pes_19_in_bits; // @[pe.scala 264:34]
  assign PE_635_io_data_0_in_valid = PENetwork_19_io_to_pes_28_in_valid; // @[pe.scala 264:34]
  assign PE_635_io_data_0_in_bits = PENetwork_19_io_to_pes_28_in_bits; // @[pe.scala 264:34]
  assign PE_636_clock = clock;
  assign PE_636_reset = reset;
  assign PE_636_io_data_2_sig_stat2trans = PENetwork_80_io_to_pes_20_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_636_io_data_1_in_valid = PENetwork_50_io_to_pes_20_in_valid; // @[pe.scala 264:34]
  assign PE_636_io_data_1_in_bits = PENetwork_50_io_to_pes_20_in_bits; // @[pe.scala 264:34]
  assign PE_636_io_data_0_in_valid = PENetwork_20_io_to_pes_28_in_valid; // @[pe.scala 264:34]
  assign PE_636_io_data_0_in_bits = PENetwork_20_io_to_pes_28_in_bits; // @[pe.scala 264:34]
  assign PE_637_clock = clock;
  assign PE_637_reset = reset;
  assign PE_637_io_data_2_sig_stat2trans = PENetwork_80_io_to_pes_21_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_637_io_data_1_in_valid = PENetwork_50_io_to_pes_21_in_valid; // @[pe.scala 264:34]
  assign PE_637_io_data_1_in_bits = PENetwork_50_io_to_pes_21_in_bits; // @[pe.scala 264:34]
  assign PE_637_io_data_0_in_valid = PENetwork_21_io_to_pes_28_in_valid; // @[pe.scala 264:34]
  assign PE_637_io_data_0_in_bits = PENetwork_21_io_to_pes_28_in_bits; // @[pe.scala 264:34]
  assign PE_638_clock = clock;
  assign PE_638_reset = reset;
  assign PE_638_io_data_2_sig_stat2trans = PENetwork_81_io_to_pes_0_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_638_io_data_1_in_valid = PENetwork_51_io_to_pes_0_in_valid; // @[pe.scala 264:34]
  assign PE_638_io_data_1_in_bits = PENetwork_51_io_to_pes_0_in_bits; // @[pe.scala 264:34]
  assign PE_638_io_data_0_in_valid = PENetwork_io_to_pes_29_in_valid; // @[pe.scala 264:34]
  assign PE_638_io_data_0_in_bits = PENetwork_io_to_pes_29_in_bits; // @[pe.scala 264:34]
  assign PE_639_clock = clock;
  assign PE_639_reset = reset;
  assign PE_639_io_data_2_sig_stat2trans = PENetwork_81_io_to_pes_1_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_639_io_data_1_in_valid = PENetwork_51_io_to_pes_1_in_valid; // @[pe.scala 264:34]
  assign PE_639_io_data_1_in_bits = PENetwork_51_io_to_pes_1_in_bits; // @[pe.scala 264:34]
  assign PE_639_io_data_0_in_valid = PENetwork_1_io_to_pes_29_in_valid; // @[pe.scala 264:34]
  assign PE_639_io_data_0_in_bits = PENetwork_1_io_to_pes_29_in_bits; // @[pe.scala 264:34]
  assign PE_640_clock = clock;
  assign PE_640_reset = reset;
  assign PE_640_io_data_2_sig_stat2trans = PENetwork_81_io_to_pes_2_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_640_io_data_1_in_valid = PENetwork_51_io_to_pes_2_in_valid; // @[pe.scala 264:34]
  assign PE_640_io_data_1_in_bits = PENetwork_51_io_to_pes_2_in_bits; // @[pe.scala 264:34]
  assign PE_640_io_data_0_in_valid = PENetwork_2_io_to_pes_29_in_valid; // @[pe.scala 264:34]
  assign PE_640_io_data_0_in_bits = PENetwork_2_io_to_pes_29_in_bits; // @[pe.scala 264:34]
  assign PE_641_clock = clock;
  assign PE_641_reset = reset;
  assign PE_641_io_data_2_sig_stat2trans = PENetwork_81_io_to_pes_3_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_641_io_data_1_in_valid = PENetwork_51_io_to_pes_3_in_valid; // @[pe.scala 264:34]
  assign PE_641_io_data_1_in_bits = PENetwork_51_io_to_pes_3_in_bits; // @[pe.scala 264:34]
  assign PE_641_io_data_0_in_valid = PENetwork_3_io_to_pes_29_in_valid; // @[pe.scala 264:34]
  assign PE_641_io_data_0_in_bits = PENetwork_3_io_to_pes_29_in_bits; // @[pe.scala 264:34]
  assign PE_642_clock = clock;
  assign PE_642_reset = reset;
  assign PE_642_io_data_2_sig_stat2trans = PENetwork_81_io_to_pes_4_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_642_io_data_1_in_valid = PENetwork_51_io_to_pes_4_in_valid; // @[pe.scala 264:34]
  assign PE_642_io_data_1_in_bits = PENetwork_51_io_to_pes_4_in_bits; // @[pe.scala 264:34]
  assign PE_642_io_data_0_in_valid = PENetwork_4_io_to_pes_29_in_valid; // @[pe.scala 264:34]
  assign PE_642_io_data_0_in_bits = PENetwork_4_io_to_pes_29_in_bits; // @[pe.scala 264:34]
  assign PE_643_clock = clock;
  assign PE_643_reset = reset;
  assign PE_643_io_data_2_sig_stat2trans = PENetwork_81_io_to_pes_5_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_643_io_data_1_in_valid = PENetwork_51_io_to_pes_5_in_valid; // @[pe.scala 264:34]
  assign PE_643_io_data_1_in_bits = PENetwork_51_io_to_pes_5_in_bits; // @[pe.scala 264:34]
  assign PE_643_io_data_0_in_valid = PENetwork_5_io_to_pes_29_in_valid; // @[pe.scala 264:34]
  assign PE_643_io_data_0_in_bits = PENetwork_5_io_to_pes_29_in_bits; // @[pe.scala 264:34]
  assign PE_644_clock = clock;
  assign PE_644_reset = reset;
  assign PE_644_io_data_2_sig_stat2trans = PENetwork_81_io_to_pes_6_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_644_io_data_1_in_valid = PENetwork_51_io_to_pes_6_in_valid; // @[pe.scala 264:34]
  assign PE_644_io_data_1_in_bits = PENetwork_51_io_to_pes_6_in_bits; // @[pe.scala 264:34]
  assign PE_644_io_data_0_in_valid = PENetwork_6_io_to_pes_29_in_valid; // @[pe.scala 264:34]
  assign PE_644_io_data_0_in_bits = PENetwork_6_io_to_pes_29_in_bits; // @[pe.scala 264:34]
  assign PE_645_clock = clock;
  assign PE_645_reset = reset;
  assign PE_645_io_data_2_sig_stat2trans = PENetwork_81_io_to_pes_7_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_645_io_data_1_in_valid = PENetwork_51_io_to_pes_7_in_valid; // @[pe.scala 264:34]
  assign PE_645_io_data_1_in_bits = PENetwork_51_io_to_pes_7_in_bits; // @[pe.scala 264:34]
  assign PE_645_io_data_0_in_valid = PENetwork_7_io_to_pes_29_in_valid; // @[pe.scala 264:34]
  assign PE_645_io_data_0_in_bits = PENetwork_7_io_to_pes_29_in_bits; // @[pe.scala 264:34]
  assign PE_646_clock = clock;
  assign PE_646_reset = reset;
  assign PE_646_io_data_2_sig_stat2trans = PENetwork_81_io_to_pes_8_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_646_io_data_1_in_valid = PENetwork_51_io_to_pes_8_in_valid; // @[pe.scala 264:34]
  assign PE_646_io_data_1_in_bits = PENetwork_51_io_to_pes_8_in_bits; // @[pe.scala 264:34]
  assign PE_646_io_data_0_in_valid = PENetwork_8_io_to_pes_29_in_valid; // @[pe.scala 264:34]
  assign PE_646_io_data_0_in_bits = PENetwork_8_io_to_pes_29_in_bits; // @[pe.scala 264:34]
  assign PE_647_clock = clock;
  assign PE_647_reset = reset;
  assign PE_647_io_data_2_sig_stat2trans = PENetwork_81_io_to_pes_9_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_647_io_data_1_in_valid = PENetwork_51_io_to_pes_9_in_valid; // @[pe.scala 264:34]
  assign PE_647_io_data_1_in_bits = PENetwork_51_io_to_pes_9_in_bits; // @[pe.scala 264:34]
  assign PE_647_io_data_0_in_valid = PENetwork_9_io_to_pes_29_in_valid; // @[pe.scala 264:34]
  assign PE_647_io_data_0_in_bits = PENetwork_9_io_to_pes_29_in_bits; // @[pe.scala 264:34]
  assign PE_648_clock = clock;
  assign PE_648_reset = reset;
  assign PE_648_io_data_2_sig_stat2trans = PENetwork_81_io_to_pes_10_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_648_io_data_1_in_valid = PENetwork_51_io_to_pes_10_in_valid; // @[pe.scala 264:34]
  assign PE_648_io_data_1_in_bits = PENetwork_51_io_to_pes_10_in_bits; // @[pe.scala 264:34]
  assign PE_648_io_data_0_in_valid = PENetwork_10_io_to_pes_29_in_valid; // @[pe.scala 264:34]
  assign PE_648_io_data_0_in_bits = PENetwork_10_io_to_pes_29_in_bits; // @[pe.scala 264:34]
  assign PE_649_clock = clock;
  assign PE_649_reset = reset;
  assign PE_649_io_data_2_sig_stat2trans = PENetwork_81_io_to_pes_11_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_649_io_data_1_in_valid = PENetwork_51_io_to_pes_11_in_valid; // @[pe.scala 264:34]
  assign PE_649_io_data_1_in_bits = PENetwork_51_io_to_pes_11_in_bits; // @[pe.scala 264:34]
  assign PE_649_io_data_0_in_valid = PENetwork_11_io_to_pes_29_in_valid; // @[pe.scala 264:34]
  assign PE_649_io_data_0_in_bits = PENetwork_11_io_to_pes_29_in_bits; // @[pe.scala 264:34]
  assign PE_650_clock = clock;
  assign PE_650_reset = reset;
  assign PE_650_io_data_2_sig_stat2trans = PENetwork_81_io_to_pes_12_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_650_io_data_1_in_valid = PENetwork_51_io_to_pes_12_in_valid; // @[pe.scala 264:34]
  assign PE_650_io_data_1_in_bits = PENetwork_51_io_to_pes_12_in_bits; // @[pe.scala 264:34]
  assign PE_650_io_data_0_in_valid = PENetwork_12_io_to_pes_29_in_valid; // @[pe.scala 264:34]
  assign PE_650_io_data_0_in_bits = PENetwork_12_io_to_pes_29_in_bits; // @[pe.scala 264:34]
  assign PE_651_clock = clock;
  assign PE_651_reset = reset;
  assign PE_651_io_data_2_sig_stat2trans = PENetwork_81_io_to_pes_13_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_651_io_data_1_in_valid = PENetwork_51_io_to_pes_13_in_valid; // @[pe.scala 264:34]
  assign PE_651_io_data_1_in_bits = PENetwork_51_io_to_pes_13_in_bits; // @[pe.scala 264:34]
  assign PE_651_io_data_0_in_valid = PENetwork_13_io_to_pes_29_in_valid; // @[pe.scala 264:34]
  assign PE_651_io_data_0_in_bits = PENetwork_13_io_to_pes_29_in_bits; // @[pe.scala 264:34]
  assign PE_652_clock = clock;
  assign PE_652_reset = reset;
  assign PE_652_io_data_2_sig_stat2trans = PENetwork_81_io_to_pes_14_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_652_io_data_1_in_valid = PENetwork_51_io_to_pes_14_in_valid; // @[pe.scala 264:34]
  assign PE_652_io_data_1_in_bits = PENetwork_51_io_to_pes_14_in_bits; // @[pe.scala 264:34]
  assign PE_652_io_data_0_in_valid = PENetwork_14_io_to_pes_29_in_valid; // @[pe.scala 264:34]
  assign PE_652_io_data_0_in_bits = PENetwork_14_io_to_pes_29_in_bits; // @[pe.scala 264:34]
  assign PE_653_clock = clock;
  assign PE_653_reset = reset;
  assign PE_653_io_data_2_sig_stat2trans = PENetwork_81_io_to_pes_15_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_653_io_data_1_in_valid = PENetwork_51_io_to_pes_15_in_valid; // @[pe.scala 264:34]
  assign PE_653_io_data_1_in_bits = PENetwork_51_io_to_pes_15_in_bits; // @[pe.scala 264:34]
  assign PE_653_io_data_0_in_valid = PENetwork_15_io_to_pes_29_in_valid; // @[pe.scala 264:34]
  assign PE_653_io_data_0_in_bits = PENetwork_15_io_to_pes_29_in_bits; // @[pe.scala 264:34]
  assign PE_654_clock = clock;
  assign PE_654_reset = reset;
  assign PE_654_io_data_2_sig_stat2trans = PENetwork_81_io_to_pes_16_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_654_io_data_1_in_valid = PENetwork_51_io_to_pes_16_in_valid; // @[pe.scala 264:34]
  assign PE_654_io_data_1_in_bits = PENetwork_51_io_to_pes_16_in_bits; // @[pe.scala 264:34]
  assign PE_654_io_data_0_in_valid = PENetwork_16_io_to_pes_29_in_valid; // @[pe.scala 264:34]
  assign PE_654_io_data_0_in_bits = PENetwork_16_io_to_pes_29_in_bits; // @[pe.scala 264:34]
  assign PE_655_clock = clock;
  assign PE_655_reset = reset;
  assign PE_655_io_data_2_sig_stat2trans = PENetwork_81_io_to_pes_17_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_655_io_data_1_in_valid = PENetwork_51_io_to_pes_17_in_valid; // @[pe.scala 264:34]
  assign PE_655_io_data_1_in_bits = PENetwork_51_io_to_pes_17_in_bits; // @[pe.scala 264:34]
  assign PE_655_io_data_0_in_valid = PENetwork_17_io_to_pes_29_in_valid; // @[pe.scala 264:34]
  assign PE_655_io_data_0_in_bits = PENetwork_17_io_to_pes_29_in_bits; // @[pe.scala 264:34]
  assign PE_656_clock = clock;
  assign PE_656_reset = reset;
  assign PE_656_io_data_2_sig_stat2trans = PENetwork_81_io_to_pes_18_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_656_io_data_1_in_valid = PENetwork_51_io_to_pes_18_in_valid; // @[pe.scala 264:34]
  assign PE_656_io_data_1_in_bits = PENetwork_51_io_to_pes_18_in_bits; // @[pe.scala 264:34]
  assign PE_656_io_data_0_in_valid = PENetwork_18_io_to_pes_29_in_valid; // @[pe.scala 264:34]
  assign PE_656_io_data_0_in_bits = PENetwork_18_io_to_pes_29_in_bits; // @[pe.scala 264:34]
  assign PE_657_clock = clock;
  assign PE_657_reset = reset;
  assign PE_657_io_data_2_sig_stat2trans = PENetwork_81_io_to_pes_19_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_657_io_data_1_in_valid = PENetwork_51_io_to_pes_19_in_valid; // @[pe.scala 264:34]
  assign PE_657_io_data_1_in_bits = PENetwork_51_io_to_pes_19_in_bits; // @[pe.scala 264:34]
  assign PE_657_io_data_0_in_valid = PENetwork_19_io_to_pes_29_in_valid; // @[pe.scala 264:34]
  assign PE_657_io_data_0_in_bits = PENetwork_19_io_to_pes_29_in_bits; // @[pe.scala 264:34]
  assign PE_658_clock = clock;
  assign PE_658_reset = reset;
  assign PE_658_io_data_2_sig_stat2trans = PENetwork_81_io_to_pes_20_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_658_io_data_1_in_valid = PENetwork_51_io_to_pes_20_in_valid; // @[pe.scala 264:34]
  assign PE_658_io_data_1_in_bits = PENetwork_51_io_to_pes_20_in_bits; // @[pe.scala 264:34]
  assign PE_658_io_data_0_in_valid = PENetwork_20_io_to_pes_29_in_valid; // @[pe.scala 264:34]
  assign PE_658_io_data_0_in_bits = PENetwork_20_io_to_pes_29_in_bits; // @[pe.scala 264:34]
  assign PE_659_clock = clock;
  assign PE_659_reset = reset;
  assign PE_659_io_data_2_sig_stat2trans = PENetwork_81_io_to_pes_21_sig_stat2trans; // @[pe.scala 266:52]
  assign PE_659_io_data_1_in_valid = PENetwork_51_io_to_pes_21_in_valid; // @[pe.scala 264:34]
  assign PE_659_io_data_1_in_bits = PENetwork_51_io_to_pes_21_in_bits; // @[pe.scala 264:34]
  assign PE_659_io_data_0_in_valid = PENetwork_21_io_to_pes_29_in_valid; // @[pe.scala 264:34]
  assign PE_659_io_data_0_in_bits = PENetwork_21_io_to_pes_29_in_bits; // @[pe.scala 264:34]
  assign PENetwork_io_to_pes_0_out_valid = PE_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_io_to_pes_0_out_bits = PE_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_io_to_pes_1_out_valid = PE_22_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_io_to_pes_1_out_bits = PE_22_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_io_to_pes_2_out_valid = PE_44_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_io_to_pes_2_out_bits = PE_44_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_io_to_pes_3_out_valid = PE_66_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_io_to_pes_3_out_bits = PE_66_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_io_to_pes_4_out_valid = PE_88_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_io_to_pes_4_out_bits = PE_88_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_io_to_pes_5_out_valid = PE_110_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_io_to_pes_5_out_bits = PE_110_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_io_to_pes_6_out_valid = PE_132_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_io_to_pes_6_out_bits = PE_132_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_io_to_pes_7_out_valid = PE_154_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_io_to_pes_7_out_bits = PE_154_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_io_to_pes_8_out_valid = PE_176_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_io_to_pes_8_out_bits = PE_176_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_io_to_pes_9_out_valid = PE_198_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_io_to_pes_9_out_bits = PE_198_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_io_to_pes_10_out_valid = PE_220_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_io_to_pes_10_out_bits = PE_220_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_io_to_pes_11_out_valid = PE_242_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_io_to_pes_11_out_bits = PE_242_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_io_to_pes_12_out_valid = PE_264_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_io_to_pes_12_out_bits = PE_264_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_io_to_pes_13_out_valid = PE_286_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_io_to_pes_13_out_bits = PE_286_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_io_to_pes_14_out_valid = PE_308_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_io_to_pes_14_out_bits = PE_308_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_io_to_pes_15_out_valid = PE_330_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_io_to_pes_15_out_bits = PE_330_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_io_to_pes_16_out_valid = PE_352_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_io_to_pes_16_out_bits = PE_352_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_io_to_pes_17_out_valid = PE_374_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_io_to_pes_17_out_bits = PE_374_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_io_to_pes_18_out_valid = PE_396_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_io_to_pes_18_out_bits = PE_396_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_io_to_pes_19_out_valid = PE_418_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_io_to_pes_19_out_bits = PE_418_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_io_to_pes_20_out_valid = PE_440_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_io_to_pes_20_out_bits = PE_440_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_io_to_pes_21_out_valid = PE_462_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_io_to_pes_21_out_bits = PE_462_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_io_to_pes_22_out_valid = PE_484_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_io_to_pes_22_out_bits = PE_484_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_io_to_pes_23_out_valid = PE_506_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_io_to_pes_23_out_bits = PE_506_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_io_to_pes_24_out_valid = PE_528_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_io_to_pes_24_out_bits = PE_528_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_io_to_pes_25_out_valid = PE_550_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_io_to_pes_25_out_bits = PE_550_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_io_to_pes_26_out_valid = PE_572_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_io_to_pes_26_out_bits = PE_572_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_io_to_pes_27_out_valid = PE_594_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_io_to_pes_27_out_bits = PE_594_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_io_to_pes_28_out_valid = PE_616_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_io_to_pes_28_out_bits = PE_616_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_io_to_mem_valid = MemController_io_rd_data_valid; // @[pe.scala 312:29]
  assign PENetwork_io_to_mem_bits = MemController_io_rd_data_bits; // @[pe.scala 312:29]
  assign PENetwork_1_io_to_pes_0_out_valid = PE_1_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_1_io_to_pes_0_out_bits = PE_1_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_1_io_to_pes_1_out_valid = PE_23_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_1_io_to_pes_1_out_bits = PE_23_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_1_io_to_pes_2_out_valid = PE_45_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_1_io_to_pes_2_out_bits = PE_45_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_1_io_to_pes_3_out_valid = PE_67_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_1_io_to_pes_3_out_bits = PE_67_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_1_io_to_pes_4_out_valid = PE_89_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_1_io_to_pes_4_out_bits = PE_89_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_1_io_to_pes_5_out_valid = PE_111_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_1_io_to_pes_5_out_bits = PE_111_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_1_io_to_pes_6_out_valid = PE_133_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_1_io_to_pes_6_out_bits = PE_133_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_1_io_to_pes_7_out_valid = PE_155_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_1_io_to_pes_7_out_bits = PE_155_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_1_io_to_pes_8_out_valid = PE_177_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_1_io_to_pes_8_out_bits = PE_177_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_1_io_to_pes_9_out_valid = PE_199_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_1_io_to_pes_9_out_bits = PE_199_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_1_io_to_pes_10_out_valid = PE_221_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_1_io_to_pes_10_out_bits = PE_221_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_1_io_to_pes_11_out_valid = PE_243_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_1_io_to_pes_11_out_bits = PE_243_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_1_io_to_pes_12_out_valid = PE_265_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_1_io_to_pes_12_out_bits = PE_265_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_1_io_to_pes_13_out_valid = PE_287_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_1_io_to_pes_13_out_bits = PE_287_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_1_io_to_pes_14_out_valid = PE_309_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_1_io_to_pes_14_out_bits = PE_309_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_1_io_to_pes_15_out_valid = PE_331_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_1_io_to_pes_15_out_bits = PE_331_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_1_io_to_pes_16_out_valid = PE_353_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_1_io_to_pes_16_out_bits = PE_353_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_1_io_to_pes_17_out_valid = PE_375_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_1_io_to_pes_17_out_bits = PE_375_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_1_io_to_pes_18_out_valid = PE_397_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_1_io_to_pes_18_out_bits = PE_397_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_1_io_to_pes_19_out_valid = PE_419_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_1_io_to_pes_19_out_bits = PE_419_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_1_io_to_pes_20_out_valid = PE_441_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_1_io_to_pes_20_out_bits = PE_441_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_1_io_to_pes_21_out_valid = PE_463_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_1_io_to_pes_21_out_bits = PE_463_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_1_io_to_pes_22_out_valid = PE_485_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_1_io_to_pes_22_out_bits = PE_485_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_1_io_to_pes_23_out_valid = PE_507_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_1_io_to_pes_23_out_bits = PE_507_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_1_io_to_pes_24_out_valid = PE_529_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_1_io_to_pes_24_out_bits = PE_529_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_1_io_to_pes_25_out_valid = PE_551_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_1_io_to_pes_25_out_bits = PE_551_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_1_io_to_pes_26_out_valid = PE_573_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_1_io_to_pes_26_out_bits = PE_573_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_1_io_to_pes_27_out_valid = PE_595_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_1_io_to_pes_27_out_bits = PE_595_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_1_io_to_pes_28_out_valid = PE_617_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_1_io_to_pes_28_out_bits = PE_617_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_1_io_to_mem_valid = MemController_1_io_rd_data_valid; // @[pe.scala 312:29]
  assign PENetwork_1_io_to_mem_bits = MemController_1_io_rd_data_bits; // @[pe.scala 312:29]
  assign PENetwork_2_io_to_pes_0_out_valid = PE_2_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_2_io_to_pes_0_out_bits = PE_2_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_2_io_to_pes_1_out_valid = PE_24_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_2_io_to_pes_1_out_bits = PE_24_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_2_io_to_pes_2_out_valid = PE_46_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_2_io_to_pes_2_out_bits = PE_46_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_2_io_to_pes_3_out_valid = PE_68_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_2_io_to_pes_3_out_bits = PE_68_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_2_io_to_pes_4_out_valid = PE_90_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_2_io_to_pes_4_out_bits = PE_90_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_2_io_to_pes_5_out_valid = PE_112_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_2_io_to_pes_5_out_bits = PE_112_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_2_io_to_pes_6_out_valid = PE_134_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_2_io_to_pes_6_out_bits = PE_134_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_2_io_to_pes_7_out_valid = PE_156_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_2_io_to_pes_7_out_bits = PE_156_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_2_io_to_pes_8_out_valid = PE_178_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_2_io_to_pes_8_out_bits = PE_178_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_2_io_to_pes_9_out_valid = PE_200_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_2_io_to_pes_9_out_bits = PE_200_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_2_io_to_pes_10_out_valid = PE_222_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_2_io_to_pes_10_out_bits = PE_222_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_2_io_to_pes_11_out_valid = PE_244_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_2_io_to_pes_11_out_bits = PE_244_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_2_io_to_pes_12_out_valid = PE_266_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_2_io_to_pes_12_out_bits = PE_266_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_2_io_to_pes_13_out_valid = PE_288_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_2_io_to_pes_13_out_bits = PE_288_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_2_io_to_pes_14_out_valid = PE_310_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_2_io_to_pes_14_out_bits = PE_310_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_2_io_to_pes_15_out_valid = PE_332_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_2_io_to_pes_15_out_bits = PE_332_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_2_io_to_pes_16_out_valid = PE_354_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_2_io_to_pes_16_out_bits = PE_354_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_2_io_to_pes_17_out_valid = PE_376_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_2_io_to_pes_17_out_bits = PE_376_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_2_io_to_pes_18_out_valid = PE_398_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_2_io_to_pes_18_out_bits = PE_398_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_2_io_to_pes_19_out_valid = PE_420_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_2_io_to_pes_19_out_bits = PE_420_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_2_io_to_pes_20_out_valid = PE_442_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_2_io_to_pes_20_out_bits = PE_442_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_2_io_to_pes_21_out_valid = PE_464_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_2_io_to_pes_21_out_bits = PE_464_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_2_io_to_pes_22_out_valid = PE_486_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_2_io_to_pes_22_out_bits = PE_486_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_2_io_to_pes_23_out_valid = PE_508_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_2_io_to_pes_23_out_bits = PE_508_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_2_io_to_pes_24_out_valid = PE_530_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_2_io_to_pes_24_out_bits = PE_530_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_2_io_to_pes_25_out_valid = PE_552_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_2_io_to_pes_25_out_bits = PE_552_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_2_io_to_pes_26_out_valid = PE_574_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_2_io_to_pes_26_out_bits = PE_574_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_2_io_to_pes_27_out_valid = PE_596_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_2_io_to_pes_27_out_bits = PE_596_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_2_io_to_pes_28_out_valid = PE_618_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_2_io_to_pes_28_out_bits = PE_618_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_2_io_to_mem_valid = MemController_2_io_rd_data_valid; // @[pe.scala 312:29]
  assign PENetwork_2_io_to_mem_bits = MemController_2_io_rd_data_bits; // @[pe.scala 312:29]
  assign PENetwork_3_io_to_pes_0_out_valid = PE_3_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_3_io_to_pes_0_out_bits = PE_3_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_3_io_to_pes_1_out_valid = PE_25_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_3_io_to_pes_1_out_bits = PE_25_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_3_io_to_pes_2_out_valid = PE_47_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_3_io_to_pes_2_out_bits = PE_47_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_3_io_to_pes_3_out_valid = PE_69_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_3_io_to_pes_3_out_bits = PE_69_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_3_io_to_pes_4_out_valid = PE_91_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_3_io_to_pes_4_out_bits = PE_91_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_3_io_to_pes_5_out_valid = PE_113_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_3_io_to_pes_5_out_bits = PE_113_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_3_io_to_pes_6_out_valid = PE_135_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_3_io_to_pes_6_out_bits = PE_135_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_3_io_to_pes_7_out_valid = PE_157_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_3_io_to_pes_7_out_bits = PE_157_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_3_io_to_pes_8_out_valid = PE_179_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_3_io_to_pes_8_out_bits = PE_179_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_3_io_to_pes_9_out_valid = PE_201_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_3_io_to_pes_9_out_bits = PE_201_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_3_io_to_pes_10_out_valid = PE_223_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_3_io_to_pes_10_out_bits = PE_223_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_3_io_to_pes_11_out_valid = PE_245_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_3_io_to_pes_11_out_bits = PE_245_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_3_io_to_pes_12_out_valid = PE_267_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_3_io_to_pes_12_out_bits = PE_267_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_3_io_to_pes_13_out_valid = PE_289_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_3_io_to_pes_13_out_bits = PE_289_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_3_io_to_pes_14_out_valid = PE_311_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_3_io_to_pes_14_out_bits = PE_311_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_3_io_to_pes_15_out_valid = PE_333_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_3_io_to_pes_15_out_bits = PE_333_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_3_io_to_pes_16_out_valid = PE_355_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_3_io_to_pes_16_out_bits = PE_355_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_3_io_to_pes_17_out_valid = PE_377_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_3_io_to_pes_17_out_bits = PE_377_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_3_io_to_pes_18_out_valid = PE_399_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_3_io_to_pes_18_out_bits = PE_399_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_3_io_to_pes_19_out_valid = PE_421_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_3_io_to_pes_19_out_bits = PE_421_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_3_io_to_pes_20_out_valid = PE_443_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_3_io_to_pes_20_out_bits = PE_443_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_3_io_to_pes_21_out_valid = PE_465_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_3_io_to_pes_21_out_bits = PE_465_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_3_io_to_pes_22_out_valid = PE_487_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_3_io_to_pes_22_out_bits = PE_487_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_3_io_to_pes_23_out_valid = PE_509_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_3_io_to_pes_23_out_bits = PE_509_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_3_io_to_pes_24_out_valid = PE_531_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_3_io_to_pes_24_out_bits = PE_531_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_3_io_to_pes_25_out_valid = PE_553_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_3_io_to_pes_25_out_bits = PE_553_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_3_io_to_pes_26_out_valid = PE_575_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_3_io_to_pes_26_out_bits = PE_575_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_3_io_to_pes_27_out_valid = PE_597_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_3_io_to_pes_27_out_bits = PE_597_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_3_io_to_pes_28_out_valid = PE_619_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_3_io_to_pes_28_out_bits = PE_619_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_3_io_to_mem_valid = MemController_3_io_rd_data_valid; // @[pe.scala 312:29]
  assign PENetwork_3_io_to_mem_bits = MemController_3_io_rd_data_bits; // @[pe.scala 312:29]
  assign PENetwork_4_io_to_pes_0_out_valid = PE_4_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_4_io_to_pes_0_out_bits = PE_4_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_4_io_to_pes_1_out_valid = PE_26_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_4_io_to_pes_1_out_bits = PE_26_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_4_io_to_pes_2_out_valid = PE_48_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_4_io_to_pes_2_out_bits = PE_48_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_4_io_to_pes_3_out_valid = PE_70_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_4_io_to_pes_3_out_bits = PE_70_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_4_io_to_pes_4_out_valid = PE_92_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_4_io_to_pes_4_out_bits = PE_92_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_4_io_to_pes_5_out_valid = PE_114_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_4_io_to_pes_5_out_bits = PE_114_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_4_io_to_pes_6_out_valid = PE_136_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_4_io_to_pes_6_out_bits = PE_136_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_4_io_to_pes_7_out_valid = PE_158_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_4_io_to_pes_7_out_bits = PE_158_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_4_io_to_pes_8_out_valid = PE_180_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_4_io_to_pes_8_out_bits = PE_180_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_4_io_to_pes_9_out_valid = PE_202_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_4_io_to_pes_9_out_bits = PE_202_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_4_io_to_pes_10_out_valid = PE_224_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_4_io_to_pes_10_out_bits = PE_224_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_4_io_to_pes_11_out_valid = PE_246_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_4_io_to_pes_11_out_bits = PE_246_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_4_io_to_pes_12_out_valid = PE_268_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_4_io_to_pes_12_out_bits = PE_268_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_4_io_to_pes_13_out_valid = PE_290_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_4_io_to_pes_13_out_bits = PE_290_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_4_io_to_pes_14_out_valid = PE_312_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_4_io_to_pes_14_out_bits = PE_312_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_4_io_to_pes_15_out_valid = PE_334_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_4_io_to_pes_15_out_bits = PE_334_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_4_io_to_pes_16_out_valid = PE_356_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_4_io_to_pes_16_out_bits = PE_356_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_4_io_to_pes_17_out_valid = PE_378_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_4_io_to_pes_17_out_bits = PE_378_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_4_io_to_pes_18_out_valid = PE_400_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_4_io_to_pes_18_out_bits = PE_400_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_4_io_to_pes_19_out_valid = PE_422_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_4_io_to_pes_19_out_bits = PE_422_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_4_io_to_pes_20_out_valid = PE_444_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_4_io_to_pes_20_out_bits = PE_444_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_4_io_to_pes_21_out_valid = PE_466_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_4_io_to_pes_21_out_bits = PE_466_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_4_io_to_pes_22_out_valid = PE_488_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_4_io_to_pes_22_out_bits = PE_488_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_4_io_to_pes_23_out_valid = PE_510_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_4_io_to_pes_23_out_bits = PE_510_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_4_io_to_pes_24_out_valid = PE_532_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_4_io_to_pes_24_out_bits = PE_532_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_4_io_to_pes_25_out_valid = PE_554_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_4_io_to_pes_25_out_bits = PE_554_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_4_io_to_pes_26_out_valid = PE_576_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_4_io_to_pes_26_out_bits = PE_576_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_4_io_to_pes_27_out_valid = PE_598_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_4_io_to_pes_27_out_bits = PE_598_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_4_io_to_pes_28_out_valid = PE_620_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_4_io_to_pes_28_out_bits = PE_620_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_4_io_to_mem_valid = MemController_4_io_rd_data_valid; // @[pe.scala 312:29]
  assign PENetwork_4_io_to_mem_bits = MemController_4_io_rd_data_bits; // @[pe.scala 312:29]
  assign PENetwork_5_io_to_pes_0_out_valid = PE_5_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_5_io_to_pes_0_out_bits = PE_5_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_5_io_to_pes_1_out_valid = PE_27_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_5_io_to_pes_1_out_bits = PE_27_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_5_io_to_pes_2_out_valid = PE_49_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_5_io_to_pes_2_out_bits = PE_49_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_5_io_to_pes_3_out_valid = PE_71_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_5_io_to_pes_3_out_bits = PE_71_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_5_io_to_pes_4_out_valid = PE_93_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_5_io_to_pes_4_out_bits = PE_93_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_5_io_to_pes_5_out_valid = PE_115_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_5_io_to_pes_5_out_bits = PE_115_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_5_io_to_pes_6_out_valid = PE_137_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_5_io_to_pes_6_out_bits = PE_137_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_5_io_to_pes_7_out_valid = PE_159_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_5_io_to_pes_7_out_bits = PE_159_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_5_io_to_pes_8_out_valid = PE_181_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_5_io_to_pes_8_out_bits = PE_181_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_5_io_to_pes_9_out_valid = PE_203_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_5_io_to_pes_9_out_bits = PE_203_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_5_io_to_pes_10_out_valid = PE_225_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_5_io_to_pes_10_out_bits = PE_225_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_5_io_to_pes_11_out_valid = PE_247_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_5_io_to_pes_11_out_bits = PE_247_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_5_io_to_pes_12_out_valid = PE_269_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_5_io_to_pes_12_out_bits = PE_269_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_5_io_to_pes_13_out_valid = PE_291_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_5_io_to_pes_13_out_bits = PE_291_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_5_io_to_pes_14_out_valid = PE_313_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_5_io_to_pes_14_out_bits = PE_313_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_5_io_to_pes_15_out_valid = PE_335_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_5_io_to_pes_15_out_bits = PE_335_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_5_io_to_pes_16_out_valid = PE_357_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_5_io_to_pes_16_out_bits = PE_357_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_5_io_to_pes_17_out_valid = PE_379_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_5_io_to_pes_17_out_bits = PE_379_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_5_io_to_pes_18_out_valid = PE_401_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_5_io_to_pes_18_out_bits = PE_401_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_5_io_to_pes_19_out_valid = PE_423_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_5_io_to_pes_19_out_bits = PE_423_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_5_io_to_pes_20_out_valid = PE_445_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_5_io_to_pes_20_out_bits = PE_445_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_5_io_to_pes_21_out_valid = PE_467_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_5_io_to_pes_21_out_bits = PE_467_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_5_io_to_pes_22_out_valid = PE_489_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_5_io_to_pes_22_out_bits = PE_489_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_5_io_to_pes_23_out_valid = PE_511_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_5_io_to_pes_23_out_bits = PE_511_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_5_io_to_pes_24_out_valid = PE_533_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_5_io_to_pes_24_out_bits = PE_533_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_5_io_to_pes_25_out_valid = PE_555_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_5_io_to_pes_25_out_bits = PE_555_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_5_io_to_pes_26_out_valid = PE_577_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_5_io_to_pes_26_out_bits = PE_577_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_5_io_to_pes_27_out_valid = PE_599_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_5_io_to_pes_27_out_bits = PE_599_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_5_io_to_pes_28_out_valid = PE_621_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_5_io_to_pes_28_out_bits = PE_621_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_5_io_to_mem_valid = MemController_5_io_rd_data_valid; // @[pe.scala 312:29]
  assign PENetwork_5_io_to_mem_bits = MemController_5_io_rd_data_bits; // @[pe.scala 312:29]
  assign PENetwork_6_io_to_pes_0_out_valid = PE_6_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_6_io_to_pes_0_out_bits = PE_6_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_6_io_to_pes_1_out_valid = PE_28_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_6_io_to_pes_1_out_bits = PE_28_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_6_io_to_pes_2_out_valid = PE_50_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_6_io_to_pes_2_out_bits = PE_50_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_6_io_to_pes_3_out_valid = PE_72_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_6_io_to_pes_3_out_bits = PE_72_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_6_io_to_pes_4_out_valid = PE_94_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_6_io_to_pes_4_out_bits = PE_94_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_6_io_to_pes_5_out_valid = PE_116_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_6_io_to_pes_5_out_bits = PE_116_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_6_io_to_pes_6_out_valid = PE_138_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_6_io_to_pes_6_out_bits = PE_138_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_6_io_to_pes_7_out_valid = PE_160_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_6_io_to_pes_7_out_bits = PE_160_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_6_io_to_pes_8_out_valid = PE_182_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_6_io_to_pes_8_out_bits = PE_182_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_6_io_to_pes_9_out_valid = PE_204_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_6_io_to_pes_9_out_bits = PE_204_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_6_io_to_pes_10_out_valid = PE_226_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_6_io_to_pes_10_out_bits = PE_226_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_6_io_to_pes_11_out_valid = PE_248_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_6_io_to_pes_11_out_bits = PE_248_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_6_io_to_pes_12_out_valid = PE_270_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_6_io_to_pes_12_out_bits = PE_270_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_6_io_to_pes_13_out_valid = PE_292_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_6_io_to_pes_13_out_bits = PE_292_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_6_io_to_pes_14_out_valid = PE_314_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_6_io_to_pes_14_out_bits = PE_314_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_6_io_to_pes_15_out_valid = PE_336_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_6_io_to_pes_15_out_bits = PE_336_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_6_io_to_pes_16_out_valid = PE_358_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_6_io_to_pes_16_out_bits = PE_358_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_6_io_to_pes_17_out_valid = PE_380_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_6_io_to_pes_17_out_bits = PE_380_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_6_io_to_pes_18_out_valid = PE_402_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_6_io_to_pes_18_out_bits = PE_402_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_6_io_to_pes_19_out_valid = PE_424_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_6_io_to_pes_19_out_bits = PE_424_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_6_io_to_pes_20_out_valid = PE_446_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_6_io_to_pes_20_out_bits = PE_446_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_6_io_to_pes_21_out_valid = PE_468_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_6_io_to_pes_21_out_bits = PE_468_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_6_io_to_pes_22_out_valid = PE_490_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_6_io_to_pes_22_out_bits = PE_490_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_6_io_to_pes_23_out_valid = PE_512_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_6_io_to_pes_23_out_bits = PE_512_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_6_io_to_pes_24_out_valid = PE_534_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_6_io_to_pes_24_out_bits = PE_534_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_6_io_to_pes_25_out_valid = PE_556_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_6_io_to_pes_25_out_bits = PE_556_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_6_io_to_pes_26_out_valid = PE_578_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_6_io_to_pes_26_out_bits = PE_578_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_6_io_to_pes_27_out_valid = PE_600_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_6_io_to_pes_27_out_bits = PE_600_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_6_io_to_pes_28_out_valid = PE_622_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_6_io_to_pes_28_out_bits = PE_622_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_6_io_to_mem_valid = MemController_6_io_rd_data_valid; // @[pe.scala 312:29]
  assign PENetwork_6_io_to_mem_bits = MemController_6_io_rd_data_bits; // @[pe.scala 312:29]
  assign PENetwork_7_io_to_pes_0_out_valid = PE_7_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_7_io_to_pes_0_out_bits = PE_7_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_7_io_to_pes_1_out_valid = PE_29_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_7_io_to_pes_1_out_bits = PE_29_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_7_io_to_pes_2_out_valid = PE_51_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_7_io_to_pes_2_out_bits = PE_51_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_7_io_to_pes_3_out_valid = PE_73_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_7_io_to_pes_3_out_bits = PE_73_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_7_io_to_pes_4_out_valid = PE_95_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_7_io_to_pes_4_out_bits = PE_95_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_7_io_to_pes_5_out_valid = PE_117_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_7_io_to_pes_5_out_bits = PE_117_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_7_io_to_pes_6_out_valid = PE_139_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_7_io_to_pes_6_out_bits = PE_139_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_7_io_to_pes_7_out_valid = PE_161_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_7_io_to_pes_7_out_bits = PE_161_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_7_io_to_pes_8_out_valid = PE_183_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_7_io_to_pes_8_out_bits = PE_183_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_7_io_to_pes_9_out_valid = PE_205_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_7_io_to_pes_9_out_bits = PE_205_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_7_io_to_pes_10_out_valid = PE_227_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_7_io_to_pes_10_out_bits = PE_227_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_7_io_to_pes_11_out_valid = PE_249_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_7_io_to_pes_11_out_bits = PE_249_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_7_io_to_pes_12_out_valid = PE_271_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_7_io_to_pes_12_out_bits = PE_271_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_7_io_to_pes_13_out_valid = PE_293_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_7_io_to_pes_13_out_bits = PE_293_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_7_io_to_pes_14_out_valid = PE_315_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_7_io_to_pes_14_out_bits = PE_315_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_7_io_to_pes_15_out_valid = PE_337_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_7_io_to_pes_15_out_bits = PE_337_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_7_io_to_pes_16_out_valid = PE_359_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_7_io_to_pes_16_out_bits = PE_359_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_7_io_to_pes_17_out_valid = PE_381_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_7_io_to_pes_17_out_bits = PE_381_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_7_io_to_pes_18_out_valid = PE_403_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_7_io_to_pes_18_out_bits = PE_403_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_7_io_to_pes_19_out_valid = PE_425_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_7_io_to_pes_19_out_bits = PE_425_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_7_io_to_pes_20_out_valid = PE_447_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_7_io_to_pes_20_out_bits = PE_447_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_7_io_to_pes_21_out_valid = PE_469_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_7_io_to_pes_21_out_bits = PE_469_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_7_io_to_pes_22_out_valid = PE_491_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_7_io_to_pes_22_out_bits = PE_491_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_7_io_to_pes_23_out_valid = PE_513_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_7_io_to_pes_23_out_bits = PE_513_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_7_io_to_pes_24_out_valid = PE_535_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_7_io_to_pes_24_out_bits = PE_535_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_7_io_to_pes_25_out_valid = PE_557_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_7_io_to_pes_25_out_bits = PE_557_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_7_io_to_pes_26_out_valid = PE_579_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_7_io_to_pes_26_out_bits = PE_579_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_7_io_to_pes_27_out_valid = PE_601_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_7_io_to_pes_27_out_bits = PE_601_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_7_io_to_pes_28_out_valid = PE_623_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_7_io_to_pes_28_out_bits = PE_623_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_7_io_to_mem_valid = MemController_7_io_rd_data_valid; // @[pe.scala 312:29]
  assign PENetwork_7_io_to_mem_bits = MemController_7_io_rd_data_bits; // @[pe.scala 312:29]
  assign PENetwork_8_io_to_pes_0_out_valid = PE_8_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_8_io_to_pes_0_out_bits = PE_8_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_8_io_to_pes_1_out_valid = PE_30_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_8_io_to_pes_1_out_bits = PE_30_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_8_io_to_pes_2_out_valid = PE_52_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_8_io_to_pes_2_out_bits = PE_52_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_8_io_to_pes_3_out_valid = PE_74_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_8_io_to_pes_3_out_bits = PE_74_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_8_io_to_pes_4_out_valid = PE_96_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_8_io_to_pes_4_out_bits = PE_96_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_8_io_to_pes_5_out_valid = PE_118_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_8_io_to_pes_5_out_bits = PE_118_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_8_io_to_pes_6_out_valid = PE_140_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_8_io_to_pes_6_out_bits = PE_140_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_8_io_to_pes_7_out_valid = PE_162_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_8_io_to_pes_7_out_bits = PE_162_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_8_io_to_pes_8_out_valid = PE_184_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_8_io_to_pes_8_out_bits = PE_184_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_8_io_to_pes_9_out_valid = PE_206_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_8_io_to_pes_9_out_bits = PE_206_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_8_io_to_pes_10_out_valid = PE_228_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_8_io_to_pes_10_out_bits = PE_228_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_8_io_to_pes_11_out_valid = PE_250_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_8_io_to_pes_11_out_bits = PE_250_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_8_io_to_pes_12_out_valid = PE_272_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_8_io_to_pes_12_out_bits = PE_272_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_8_io_to_pes_13_out_valid = PE_294_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_8_io_to_pes_13_out_bits = PE_294_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_8_io_to_pes_14_out_valid = PE_316_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_8_io_to_pes_14_out_bits = PE_316_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_8_io_to_pes_15_out_valid = PE_338_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_8_io_to_pes_15_out_bits = PE_338_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_8_io_to_pes_16_out_valid = PE_360_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_8_io_to_pes_16_out_bits = PE_360_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_8_io_to_pes_17_out_valid = PE_382_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_8_io_to_pes_17_out_bits = PE_382_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_8_io_to_pes_18_out_valid = PE_404_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_8_io_to_pes_18_out_bits = PE_404_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_8_io_to_pes_19_out_valid = PE_426_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_8_io_to_pes_19_out_bits = PE_426_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_8_io_to_pes_20_out_valid = PE_448_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_8_io_to_pes_20_out_bits = PE_448_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_8_io_to_pes_21_out_valid = PE_470_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_8_io_to_pes_21_out_bits = PE_470_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_8_io_to_pes_22_out_valid = PE_492_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_8_io_to_pes_22_out_bits = PE_492_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_8_io_to_pes_23_out_valid = PE_514_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_8_io_to_pes_23_out_bits = PE_514_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_8_io_to_pes_24_out_valid = PE_536_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_8_io_to_pes_24_out_bits = PE_536_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_8_io_to_pes_25_out_valid = PE_558_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_8_io_to_pes_25_out_bits = PE_558_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_8_io_to_pes_26_out_valid = PE_580_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_8_io_to_pes_26_out_bits = PE_580_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_8_io_to_pes_27_out_valid = PE_602_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_8_io_to_pes_27_out_bits = PE_602_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_8_io_to_pes_28_out_valid = PE_624_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_8_io_to_pes_28_out_bits = PE_624_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_8_io_to_mem_valid = MemController_8_io_rd_data_valid; // @[pe.scala 312:29]
  assign PENetwork_8_io_to_mem_bits = MemController_8_io_rd_data_bits; // @[pe.scala 312:29]
  assign PENetwork_9_io_to_pes_0_out_valid = PE_9_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_9_io_to_pes_0_out_bits = PE_9_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_9_io_to_pes_1_out_valid = PE_31_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_9_io_to_pes_1_out_bits = PE_31_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_9_io_to_pes_2_out_valid = PE_53_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_9_io_to_pes_2_out_bits = PE_53_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_9_io_to_pes_3_out_valid = PE_75_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_9_io_to_pes_3_out_bits = PE_75_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_9_io_to_pes_4_out_valid = PE_97_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_9_io_to_pes_4_out_bits = PE_97_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_9_io_to_pes_5_out_valid = PE_119_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_9_io_to_pes_5_out_bits = PE_119_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_9_io_to_pes_6_out_valid = PE_141_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_9_io_to_pes_6_out_bits = PE_141_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_9_io_to_pes_7_out_valid = PE_163_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_9_io_to_pes_7_out_bits = PE_163_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_9_io_to_pes_8_out_valid = PE_185_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_9_io_to_pes_8_out_bits = PE_185_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_9_io_to_pes_9_out_valid = PE_207_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_9_io_to_pes_9_out_bits = PE_207_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_9_io_to_pes_10_out_valid = PE_229_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_9_io_to_pes_10_out_bits = PE_229_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_9_io_to_pes_11_out_valid = PE_251_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_9_io_to_pes_11_out_bits = PE_251_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_9_io_to_pes_12_out_valid = PE_273_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_9_io_to_pes_12_out_bits = PE_273_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_9_io_to_pes_13_out_valid = PE_295_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_9_io_to_pes_13_out_bits = PE_295_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_9_io_to_pes_14_out_valid = PE_317_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_9_io_to_pes_14_out_bits = PE_317_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_9_io_to_pes_15_out_valid = PE_339_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_9_io_to_pes_15_out_bits = PE_339_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_9_io_to_pes_16_out_valid = PE_361_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_9_io_to_pes_16_out_bits = PE_361_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_9_io_to_pes_17_out_valid = PE_383_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_9_io_to_pes_17_out_bits = PE_383_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_9_io_to_pes_18_out_valid = PE_405_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_9_io_to_pes_18_out_bits = PE_405_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_9_io_to_pes_19_out_valid = PE_427_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_9_io_to_pes_19_out_bits = PE_427_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_9_io_to_pes_20_out_valid = PE_449_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_9_io_to_pes_20_out_bits = PE_449_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_9_io_to_pes_21_out_valid = PE_471_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_9_io_to_pes_21_out_bits = PE_471_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_9_io_to_pes_22_out_valid = PE_493_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_9_io_to_pes_22_out_bits = PE_493_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_9_io_to_pes_23_out_valid = PE_515_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_9_io_to_pes_23_out_bits = PE_515_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_9_io_to_pes_24_out_valid = PE_537_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_9_io_to_pes_24_out_bits = PE_537_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_9_io_to_pes_25_out_valid = PE_559_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_9_io_to_pes_25_out_bits = PE_559_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_9_io_to_pes_26_out_valid = PE_581_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_9_io_to_pes_26_out_bits = PE_581_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_9_io_to_pes_27_out_valid = PE_603_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_9_io_to_pes_27_out_bits = PE_603_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_9_io_to_pes_28_out_valid = PE_625_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_9_io_to_pes_28_out_bits = PE_625_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_9_io_to_mem_valid = MemController_9_io_rd_data_valid; // @[pe.scala 312:29]
  assign PENetwork_9_io_to_mem_bits = MemController_9_io_rd_data_bits; // @[pe.scala 312:29]
  assign PENetwork_10_io_to_pes_0_out_valid = PE_10_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_10_io_to_pes_0_out_bits = PE_10_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_10_io_to_pes_1_out_valid = PE_32_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_10_io_to_pes_1_out_bits = PE_32_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_10_io_to_pes_2_out_valid = PE_54_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_10_io_to_pes_2_out_bits = PE_54_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_10_io_to_pes_3_out_valid = PE_76_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_10_io_to_pes_3_out_bits = PE_76_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_10_io_to_pes_4_out_valid = PE_98_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_10_io_to_pes_4_out_bits = PE_98_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_10_io_to_pes_5_out_valid = PE_120_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_10_io_to_pes_5_out_bits = PE_120_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_10_io_to_pes_6_out_valid = PE_142_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_10_io_to_pes_6_out_bits = PE_142_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_10_io_to_pes_7_out_valid = PE_164_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_10_io_to_pes_7_out_bits = PE_164_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_10_io_to_pes_8_out_valid = PE_186_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_10_io_to_pes_8_out_bits = PE_186_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_10_io_to_pes_9_out_valid = PE_208_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_10_io_to_pes_9_out_bits = PE_208_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_10_io_to_pes_10_out_valid = PE_230_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_10_io_to_pes_10_out_bits = PE_230_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_10_io_to_pes_11_out_valid = PE_252_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_10_io_to_pes_11_out_bits = PE_252_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_10_io_to_pes_12_out_valid = PE_274_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_10_io_to_pes_12_out_bits = PE_274_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_10_io_to_pes_13_out_valid = PE_296_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_10_io_to_pes_13_out_bits = PE_296_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_10_io_to_pes_14_out_valid = PE_318_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_10_io_to_pes_14_out_bits = PE_318_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_10_io_to_pes_15_out_valid = PE_340_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_10_io_to_pes_15_out_bits = PE_340_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_10_io_to_pes_16_out_valid = PE_362_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_10_io_to_pes_16_out_bits = PE_362_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_10_io_to_pes_17_out_valid = PE_384_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_10_io_to_pes_17_out_bits = PE_384_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_10_io_to_pes_18_out_valid = PE_406_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_10_io_to_pes_18_out_bits = PE_406_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_10_io_to_pes_19_out_valid = PE_428_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_10_io_to_pes_19_out_bits = PE_428_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_10_io_to_pes_20_out_valid = PE_450_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_10_io_to_pes_20_out_bits = PE_450_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_10_io_to_pes_21_out_valid = PE_472_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_10_io_to_pes_21_out_bits = PE_472_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_10_io_to_pes_22_out_valid = PE_494_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_10_io_to_pes_22_out_bits = PE_494_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_10_io_to_pes_23_out_valid = PE_516_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_10_io_to_pes_23_out_bits = PE_516_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_10_io_to_pes_24_out_valid = PE_538_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_10_io_to_pes_24_out_bits = PE_538_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_10_io_to_pes_25_out_valid = PE_560_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_10_io_to_pes_25_out_bits = PE_560_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_10_io_to_pes_26_out_valid = PE_582_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_10_io_to_pes_26_out_bits = PE_582_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_10_io_to_pes_27_out_valid = PE_604_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_10_io_to_pes_27_out_bits = PE_604_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_10_io_to_pes_28_out_valid = PE_626_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_10_io_to_pes_28_out_bits = PE_626_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_10_io_to_mem_valid = MemController_10_io_rd_data_valid; // @[pe.scala 312:29]
  assign PENetwork_10_io_to_mem_bits = MemController_10_io_rd_data_bits; // @[pe.scala 312:29]
  assign PENetwork_11_io_to_pes_0_out_valid = PE_11_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_11_io_to_pes_0_out_bits = PE_11_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_11_io_to_pes_1_out_valid = PE_33_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_11_io_to_pes_1_out_bits = PE_33_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_11_io_to_pes_2_out_valid = PE_55_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_11_io_to_pes_2_out_bits = PE_55_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_11_io_to_pes_3_out_valid = PE_77_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_11_io_to_pes_3_out_bits = PE_77_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_11_io_to_pes_4_out_valid = PE_99_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_11_io_to_pes_4_out_bits = PE_99_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_11_io_to_pes_5_out_valid = PE_121_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_11_io_to_pes_5_out_bits = PE_121_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_11_io_to_pes_6_out_valid = PE_143_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_11_io_to_pes_6_out_bits = PE_143_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_11_io_to_pes_7_out_valid = PE_165_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_11_io_to_pes_7_out_bits = PE_165_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_11_io_to_pes_8_out_valid = PE_187_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_11_io_to_pes_8_out_bits = PE_187_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_11_io_to_pes_9_out_valid = PE_209_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_11_io_to_pes_9_out_bits = PE_209_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_11_io_to_pes_10_out_valid = PE_231_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_11_io_to_pes_10_out_bits = PE_231_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_11_io_to_pes_11_out_valid = PE_253_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_11_io_to_pes_11_out_bits = PE_253_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_11_io_to_pes_12_out_valid = PE_275_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_11_io_to_pes_12_out_bits = PE_275_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_11_io_to_pes_13_out_valid = PE_297_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_11_io_to_pes_13_out_bits = PE_297_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_11_io_to_pes_14_out_valid = PE_319_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_11_io_to_pes_14_out_bits = PE_319_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_11_io_to_pes_15_out_valid = PE_341_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_11_io_to_pes_15_out_bits = PE_341_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_11_io_to_pes_16_out_valid = PE_363_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_11_io_to_pes_16_out_bits = PE_363_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_11_io_to_pes_17_out_valid = PE_385_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_11_io_to_pes_17_out_bits = PE_385_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_11_io_to_pes_18_out_valid = PE_407_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_11_io_to_pes_18_out_bits = PE_407_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_11_io_to_pes_19_out_valid = PE_429_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_11_io_to_pes_19_out_bits = PE_429_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_11_io_to_pes_20_out_valid = PE_451_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_11_io_to_pes_20_out_bits = PE_451_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_11_io_to_pes_21_out_valid = PE_473_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_11_io_to_pes_21_out_bits = PE_473_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_11_io_to_pes_22_out_valid = PE_495_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_11_io_to_pes_22_out_bits = PE_495_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_11_io_to_pes_23_out_valid = PE_517_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_11_io_to_pes_23_out_bits = PE_517_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_11_io_to_pes_24_out_valid = PE_539_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_11_io_to_pes_24_out_bits = PE_539_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_11_io_to_pes_25_out_valid = PE_561_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_11_io_to_pes_25_out_bits = PE_561_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_11_io_to_pes_26_out_valid = PE_583_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_11_io_to_pes_26_out_bits = PE_583_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_11_io_to_pes_27_out_valid = PE_605_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_11_io_to_pes_27_out_bits = PE_605_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_11_io_to_pes_28_out_valid = PE_627_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_11_io_to_pes_28_out_bits = PE_627_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_11_io_to_mem_valid = MemController_11_io_rd_data_valid; // @[pe.scala 312:29]
  assign PENetwork_11_io_to_mem_bits = MemController_11_io_rd_data_bits; // @[pe.scala 312:29]
  assign PENetwork_12_io_to_pes_0_out_valid = PE_12_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_12_io_to_pes_0_out_bits = PE_12_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_12_io_to_pes_1_out_valid = PE_34_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_12_io_to_pes_1_out_bits = PE_34_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_12_io_to_pes_2_out_valid = PE_56_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_12_io_to_pes_2_out_bits = PE_56_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_12_io_to_pes_3_out_valid = PE_78_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_12_io_to_pes_3_out_bits = PE_78_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_12_io_to_pes_4_out_valid = PE_100_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_12_io_to_pes_4_out_bits = PE_100_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_12_io_to_pes_5_out_valid = PE_122_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_12_io_to_pes_5_out_bits = PE_122_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_12_io_to_pes_6_out_valid = PE_144_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_12_io_to_pes_6_out_bits = PE_144_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_12_io_to_pes_7_out_valid = PE_166_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_12_io_to_pes_7_out_bits = PE_166_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_12_io_to_pes_8_out_valid = PE_188_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_12_io_to_pes_8_out_bits = PE_188_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_12_io_to_pes_9_out_valid = PE_210_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_12_io_to_pes_9_out_bits = PE_210_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_12_io_to_pes_10_out_valid = PE_232_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_12_io_to_pes_10_out_bits = PE_232_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_12_io_to_pes_11_out_valid = PE_254_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_12_io_to_pes_11_out_bits = PE_254_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_12_io_to_pes_12_out_valid = PE_276_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_12_io_to_pes_12_out_bits = PE_276_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_12_io_to_pes_13_out_valid = PE_298_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_12_io_to_pes_13_out_bits = PE_298_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_12_io_to_pes_14_out_valid = PE_320_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_12_io_to_pes_14_out_bits = PE_320_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_12_io_to_pes_15_out_valid = PE_342_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_12_io_to_pes_15_out_bits = PE_342_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_12_io_to_pes_16_out_valid = PE_364_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_12_io_to_pes_16_out_bits = PE_364_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_12_io_to_pes_17_out_valid = PE_386_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_12_io_to_pes_17_out_bits = PE_386_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_12_io_to_pes_18_out_valid = PE_408_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_12_io_to_pes_18_out_bits = PE_408_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_12_io_to_pes_19_out_valid = PE_430_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_12_io_to_pes_19_out_bits = PE_430_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_12_io_to_pes_20_out_valid = PE_452_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_12_io_to_pes_20_out_bits = PE_452_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_12_io_to_pes_21_out_valid = PE_474_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_12_io_to_pes_21_out_bits = PE_474_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_12_io_to_pes_22_out_valid = PE_496_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_12_io_to_pes_22_out_bits = PE_496_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_12_io_to_pes_23_out_valid = PE_518_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_12_io_to_pes_23_out_bits = PE_518_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_12_io_to_pes_24_out_valid = PE_540_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_12_io_to_pes_24_out_bits = PE_540_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_12_io_to_pes_25_out_valid = PE_562_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_12_io_to_pes_25_out_bits = PE_562_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_12_io_to_pes_26_out_valid = PE_584_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_12_io_to_pes_26_out_bits = PE_584_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_12_io_to_pes_27_out_valid = PE_606_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_12_io_to_pes_27_out_bits = PE_606_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_12_io_to_pes_28_out_valid = PE_628_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_12_io_to_pes_28_out_bits = PE_628_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_12_io_to_mem_valid = MemController_12_io_rd_data_valid; // @[pe.scala 312:29]
  assign PENetwork_12_io_to_mem_bits = MemController_12_io_rd_data_bits; // @[pe.scala 312:29]
  assign PENetwork_13_io_to_pes_0_out_valid = PE_13_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_13_io_to_pes_0_out_bits = PE_13_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_13_io_to_pes_1_out_valid = PE_35_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_13_io_to_pes_1_out_bits = PE_35_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_13_io_to_pes_2_out_valid = PE_57_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_13_io_to_pes_2_out_bits = PE_57_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_13_io_to_pes_3_out_valid = PE_79_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_13_io_to_pes_3_out_bits = PE_79_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_13_io_to_pes_4_out_valid = PE_101_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_13_io_to_pes_4_out_bits = PE_101_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_13_io_to_pes_5_out_valid = PE_123_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_13_io_to_pes_5_out_bits = PE_123_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_13_io_to_pes_6_out_valid = PE_145_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_13_io_to_pes_6_out_bits = PE_145_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_13_io_to_pes_7_out_valid = PE_167_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_13_io_to_pes_7_out_bits = PE_167_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_13_io_to_pes_8_out_valid = PE_189_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_13_io_to_pes_8_out_bits = PE_189_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_13_io_to_pes_9_out_valid = PE_211_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_13_io_to_pes_9_out_bits = PE_211_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_13_io_to_pes_10_out_valid = PE_233_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_13_io_to_pes_10_out_bits = PE_233_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_13_io_to_pes_11_out_valid = PE_255_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_13_io_to_pes_11_out_bits = PE_255_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_13_io_to_pes_12_out_valid = PE_277_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_13_io_to_pes_12_out_bits = PE_277_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_13_io_to_pes_13_out_valid = PE_299_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_13_io_to_pes_13_out_bits = PE_299_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_13_io_to_pes_14_out_valid = PE_321_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_13_io_to_pes_14_out_bits = PE_321_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_13_io_to_pes_15_out_valid = PE_343_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_13_io_to_pes_15_out_bits = PE_343_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_13_io_to_pes_16_out_valid = PE_365_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_13_io_to_pes_16_out_bits = PE_365_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_13_io_to_pes_17_out_valid = PE_387_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_13_io_to_pes_17_out_bits = PE_387_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_13_io_to_pes_18_out_valid = PE_409_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_13_io_to_pes_18_out_bits = PE_409_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_13_io_to_pes_19_out_valid = PE_431_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_13_io_to_pes_19_out_bits = PE_431_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_13_io_to_pes_20_out_valid = PE_453_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_13_io_to_pes_20_out_bits = PE_453_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_13_io_to_pes_21_out_valid = PE_475_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_13_io_to_pes_21_out_bits = PE_475_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_13_io_to_pes_22_out_valid = PE_497_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_13_io_to_pes_22_out_bits = PE_497_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_13_io_to_pes_23_out_valid = PE_519_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_13_io_to_pes_23_out_bits = PE_519_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_13_io_to_pes_24_out_valid = PE_541_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_13_io_to_pes_24_out_bits = PE_541_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_13_io_to_pes_25_out_valid = PE_563_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_13_io_to_pes_25_out_bits = PE_563_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_13_io_to_pes_26_out_valid = PE_585_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_13_io_to_pes_26_out_bits = PE_585_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_13_io_to_pes_27_out_valid = PE_607_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_13_io_to_pes_27_out_bits = PE_607_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_13_io_to_pes_28_out_valid = PE_629_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_13_io_to_pes_28_out_bits = PE_629_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_13_io_to_mem_valid = MemController_13_io_rd_data_valid; // @[pe.scala 312:29]
  assign PENetwork_13_io_to_mem_bits = MemController_13_io_rd_data_bits; // @[pe.scala 312:29]
  assign PENetwork_14_io_to_pes_0_out_valid = PE_14_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_14_io_to_pes_0_out_bits = PE_14_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_14_io_to_pes_1_out_valid = PE_36_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_14_io_to_pes_1_out_bits = PE_36_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_14_io_to_pes_2_out_valid = PE_58_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_14_io_to_pes_2_out_bits = PE_58_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_14_io_to_pes_3_out_valid = PE_80_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_14_io_to_pes_3_out_bits = PE_80_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_14_io_to_pes_4_out_valid = PE_102_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_14_io_to_pes_4_out_bits = PE_102_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_14_io_to_pes_5_out_valid = PE_124_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_14_io_to_pes_5_out_bits = PE_124_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_14_io_to_pes_6_out_valid = PE_146_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_14_io_to_pes_6_out_bits = PE_146_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_14_io_to_pes_7_out_valid = PE_168_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_14_io_to_pes_7_out_bits = PE_168_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_14_io_to_pes_8_out_valid = PE_190_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_14_io_to_pes_8_out_bits = PE_190_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_14_io_to_pes_9_out_valid = PE_212_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_14_io_to_pes_9_out_bits = PE_212_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_14_io_to_pes_10_out_valid = PE_234_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_14_io_to_pes_10_out_bits = PE_234_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_14_io_to_pes_11_out_valid = PE_256_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_14_io_to_pes_11_out_bits = PE_256_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_14_io_to_pes_12_out_valid = PE_278_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_14_io_to_pes_12_out_bits = PE_278_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_14_io_to_pes_13_out_valid = PE_300_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_14_io_to_pes_13_out_bits = PE_300_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_14_io_to_pes_14_out_valid = PE_322_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_14_io_to_pes_14_out_bits = PE_322_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_14_io_to_pes_15_out_valid = PE_344_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_14_io_to_pes_15_out_bits = PE_344_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_14_io_to_pes_16_out_valid = PE_366_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_14_io_to_pes_16_out_bits = PE_366_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_14_io_to_pes_17_out_valid = PE_388_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_14_io_to_pes_17_out_bits = PE_388_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_14_io_to_pes_18_out_valid = PE_410_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_14_io_to_pes_18_out_bits = PE_410_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_14_io_to_pes_19_out_valid = PE_432_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_14_io_to_pes_19_out_bits = PE_432_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_14_io_to_pes_20_out_valid = PE_454_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_14_io_to_pes_20_out_bits = PE_454_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_14_io_to_pes_21_out_valid = PE_476_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_14_io_to_pes_21_out_bits = PE_476_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_14_io_to_pes_22_out_valid = PE_498_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_14_io_to_pes_22_out_bits = PE_498_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_14_io_to_pes_23_out_valid = PE_520_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_14_io_to_pes_23_out_bits = PE_520_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_14_io_to_pes_24_out_valid = PE_542_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_14_io_to_pes_24_out_bits = PE_542_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_14_io_to_pes_25_out_valid = PE_564_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_14_io_to_pes_25_out_bits = PE_564_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_14_io_to_pes_26_out_valid = PE_586_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_14_io_to_pes_26_out_bits = PE_586_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_14_io_to_pes_27_out_valid = PE_608_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_14_io_to_pes_27_out_bits = PE_608_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_14_io_to_pes_28_out_valid = PE_630_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_14_io_to_pes_28_out_bits = PE_630_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_14_io_to_mem_valid = MemController_14_io_rd_data_valid; // @[pe.scala 312:29]
  assign PENetwork_14_io_to_mem_bits = MemController_14_io_rd_data_bits; // @[pe.scala 312:29]
  assign PENetwork_15_io_to_pes_0_out_valid = PE_15_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_15_io_to_pes_0_out_bits = PE_15_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_15_io_to_pes_1_out_valid = PE_37_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_15_io_to_pes_1_out_bits = PE_37_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_15_io_to_pes_2_out_valid = PE_59_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_15_io_to_pes_2_out_bits = PE_59_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_15_io_to_pes_3_out_valid = PE_81_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_15_io_to_pes_3_out_bits = PE_81_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_15_io_to_pes_4_out_valid = PE_103_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_15_io_to_pes_4_out_bits = PE_103_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_15_io_to_pes_5_out_valid = PE_125_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_15_io_to_pes_5_out_bits = PE_125_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_15_io_to_pes_6_out_valid = PE_147_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_15_io_to_pes_6_out_bits = PE_147_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_15_io_to_pes_7_out_valid = PE_169_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_15_io_to_pes_7_out_bits = PE_169_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_15_io_to_pes_8_out_valid = PE_191_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_15_io_to_pes_8_out_bits = PE_191_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_15_io_to_pes_9_out_valid = PE_213_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_15_io_to_pes_9_out_bits = PE_213_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_15_io_to_pes_10_out_valid = PE_235_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_15_io_to_pes_10_out_bits = PE_235_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_15_io_to_pes_11_out_valid = PE_257_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_15_io_to_pes_11_out_bits = PE_257_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_15_io_to_pes_12_out_valid = PE_279_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_15_io_to_pes_12_out_bits = PE_279_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_15_io_to_pes_13_out_valid = PE_301_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_15_io_to_pes_13_out_bits = PE_301_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_15_io_to_pes_14_out_valid = PE_323_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_15_io_to_pes_14_out_bits = PE_323_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_15_io_to_pes_15_out_valid = PE_345_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_15_io_to_pes_15_out_bits = PE_345_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_15_io_to_pes_16_out_valid = PE_367_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_15_io_to_pes_16_out_bits = PE_367_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_15_io_to_pes_17_out_valid = PE_389_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_15_io_to_pes_17_out_bits = PE_389_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_15_io_to_pes_18_out_valid = PE_411_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_15_io_to_pes_18_out_bits = PE_411_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_15_io_to_pes_19_out_valid = PE_433_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_15_io_to_pes_19_out_bits = PE_433_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_15_io_to_pes_20_out_valid = PE_455_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_15_io_to_pes_20_out_bits = PE_455_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_15_io_to_pes_21_out_valid = PE_477_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_15_io_to_pes_21_out_bits = PE_477_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_15_io_to_pes_22_out_valid = PE_499_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_15_io_to_pes_22_out_bits = PE_499_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_15_io_to_pes_23_out_valid = PE_521_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_15_io_to_pes_23_out_bits = PE_521_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_15_io_to_pes_24_out_valid = PE_543_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_15_io_to_pes_24_out_bits = PE_543_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_15_io_to_pes_25_out_valid = PE_565_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_15_io_to_pes_25_out_bits = PE_565_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_15_io_to_pes_26_out_valid = PE_587_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_15_io_to_pes_26_out_bits = PE_587_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_15_io_to_pes_27_out_valid = PE_609_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_15_io_to_pes_27_out_bits = PE_609_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_15_io_to_pes_28_out_valid = PE_631_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_15_io_to_pes_28_out_bits = PE_631_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_15_io_to_mem_valid = MemController_15_io_rd_data_valid; // @[pe.scala 312:29]
  assign PENetwork_15_io_to_mem_bits = MemController_15_io_rd_data_bits; // @[pe.scala 312:29]
  assign PENetwork_16_io_to_pes_0_out_valid = PE_16_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_16_io_to_pes_0_out_bits = PE_16_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_16_io_to_pes_1_out_valid = PE_38_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_16_io_to_pes_1_out_bits = PE_38_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_16_io_to_pes_2_out_valid = PE_60_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_16_io_to_pes_2_out_bits = PE_60_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_16_io_to_pes_3_out_valid = PE_82_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_16_io_to_pes_3_out_bits = PE_82_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_16_io_to_pes_4_out_valid = PE_104_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_16_io_to_pes_4_out_bits = PE_104_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_16_io_to_pes_5_out_valid = PE_126_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_16_io_to_pes_5_out_bits = PE_126_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_16_io_to_pes_6_out_valid = PE_148_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_16_io_to_pes_6_out_bits = PE_148_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_16_io_to_pes_7_out_valid = PE_170_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_16_io_to_pes_7_out_bits = PE_170_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_16_io_to_pes_8_out_valid = PE_192_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_16_io_to_pes_8_out_bits = PE_192_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_16_io_to_pes_9_out_valid = PE_214_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_16_io_to_pes_9_out_bits = PE_214_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_16_io_to_pes_10_out_valid = PE_236_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_16_io_to_pes_10_out_bits = PE_236_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_16_io_to_pes_11_out_valid = PE_258_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_16_io_to_pes_11_out_bits = PE_258_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_16_io_to_pes_12_out_valid = PE_280_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_16_io_to_pes_12_out_bits = PE_280_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_16_io_to_pes_13_out_valid = PE_302_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_16_io_to_pes_13_out_bits = PE_302_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_16_io_to_pes_14_out_valid = PE_324_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_16_io_to_pes_14_out_bits = PE_324_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_16_io_to_pes_15_out_valid = PE_346_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_16_io_to_pes_15_out_bits = PE_346_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_16_io_to_pes_16_out_valid = PE_368_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_16_io_to_pes_16_out_bits = PE_368_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_16_io_to_pes_17_out_valid = PE_390_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_16_io_to_pes_17_out_bits = PE_390_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_16_io_to_pes_18_out_valid = PE_412_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_16_io_to_pes_18_out_bits = PE_412_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_16_io_to_pes_19_out_valid = PE_434_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_16_io_to_pes_19_out_bits = PE_434_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_16_io_to_pes_20_out_valid = PE_456_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_16_io_to_pes_20_out_bits = PE_456_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_16_io_to_pes_21_out_valid = PE_478_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_16_io_to_pes_21_out_bits = PE_478_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_16_io_to_pes_22_out_valid = PE_500_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_16_io_to_pes_22_out_bits = PE_500_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_16_io_to_pes_23_out_valid = PE_522_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_16_io_to_pes_23_out_bits = PE_522_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_16_io_to_pes_24_out_valid = PE_544_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_16_io_to_pes_24_out_bits = PE_544_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_16_io_to_pes_25_out_valid = PE_566_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_16_io_to_pes_25_out_bits = PE_566_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_16_io_to_pes_26_out_valid = PE_588_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_16_io_to_pes_26_out_bits = PE_588_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_16_io_to_pes_27_out_valid = PE_610_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_16_io_to_pes_27_out_bits = PE_610_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_16_io_to_pes_28_out_valid = PE_632_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_16_io_to_pes_28_out_bits = PE_632_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_16_io_to_mem_valid = MemController_16_io_rd_data_valid; // @[pe.scala 312:29]
  assign PENetwork_16_io_to_mem_bits = MemController_16_io_rd_data_bits; // @[pe.scala 312:29]
  assign PENetwork_17_io_to_pes_0_out_valid = PE_17_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_17_io_to_pes_0_out_bits = PE_17_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_17_io_to_pes_1_out_valid = PE_39_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_17_io_to_pes_1_out_bits = PE_39_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_17_io_to_pes_2_out_valid = PE_61_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_17_io_to_pes_2_out_bits = PE_61_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_17_io_to_pes_3_out_valid = PE_83_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_17_io_to_pes_3_out_bits = PE_83_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_17_io_to_pes_4_out_valid = PE_105_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_17_io_to_pes_4_out_bits = PE_105_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_17_io_to_pes_5_out_valid = PE_127_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_17_io_to_pes_5_out_bits = PE_127_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_17_io_to_pes_6_out_valid = PE_149_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_17_io_to_pes_6_out_bits = PE_149_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_17_io_to_pes_7_out_valid = PE_171_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_17_io_to_pes_7_out_bits = PE_171_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_17_io_to_pes_8_out_valid = PE_193_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_17_io_to_pes_8_out_bits = PE_193_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_17_io_to_pes_9_out_valid = PE_215_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_17_io_to_pes_9_out_bits = PE_215_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_17_io_to_pes_10_out_valid = PE_237_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_17_io_to_pes_10_out_bits = PE_237_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_17_io_to_pes_11_out_valid = PE_259_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_17_io_to_pes_11_out_bits = PE_259_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_17_io_to_pes_12_out_valid = PE_281_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_17_io_to_pes_12_out_bits = PE_281_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_17_io_to_pes_13_out_valid = PE_303_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_17_io_to_pes_13_out_bits = PE_303_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_17_io_to_pes_14_out_valid = PE_325_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_17_io_to_pes_14_out_bits = PE_325_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_17_io_to_pes_15_out_valid = PE_347_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_17_io_to_pes_15_out_bits = PE_347_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_17_io_to_pes_16_out_valid = PE_369_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_17_io_to_pes_16_out_bits = PE_369_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_17_io_to_pes_17_out_valid = PE_391_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_17_io_to_pes_17_out_bits = PE_391_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_17_io_to_pes_18_out_valid = PE_413_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_17_io_to_pes_18_out_bits = PE_413_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_17_io_to_pes_19_out_valid = PE_435_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_17_io_to_pes_19_out_bits = PE_435_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_17_io_to_pes_20_out_valid = PE_457_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_17_io_to_pes_20_out_bits = PE_457_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_17_io_to_pes_21_out_valid = PE_479_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_17_io_to_pes_21_out_bits = PE_479_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_17_io_to_pes_22_out_valid = PE_501_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_17_io_to_pes_22_out_bits = PE_501_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_17_io_to_pes_23_out_valid = PE_523_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_17_io_to_pes_23_out_bits = PE_523_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_17_io_to_pes_24_out_valid = PE_545_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_17_io_to_pes_24_out_bits = PE_545_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_17_io_to_pes_25_out_valid = PE_567_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_17_io_to_pes_25_out_bits = PE_567_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_17_io_to_pes_26_out_valid = PE_589_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_17_io_to_pes_26_out_bits = PE_589_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_17_io_to_pes_27_out_valid = PE_611_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_17_io_to_pes_27_out_bits = PE_611_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_17_io_to_pes_28_out_valid = PE_633_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_17_io_to_pes_28_out_bits = PE_633_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_17_io_to_mem_valid = MemController_17_io_rd_data_valid; // @[pe.scala 312:29]
  assign PENetwork_17_io_to_mem_bits = MemController_17_io_rd_data_bits; // @[pe.scala 312:29]
  assign PENetwork_18_io_to_pes_0_out_valid = PE_18_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_18_io_to_pes_0_out_bits = PE_18_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_18_io_to_pes_1_out_valid = PE_40_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_18_io_to_pes_1_out_bits = PE_40_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_18_io_to_pes_2_out_valid = PE_62_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_18_io_to_pes_2_out_bits = PE_62_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_18_io_to_pes_3_out_valid = PE_84_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_18_io_to_pes_3_out_bits = PE_84_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_18_io_to_pes_4_out_valid = PE_106_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_18_io_to_pes_4_out_bits = PE_106_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_18_io_to_pes_5_out_valid = PE_128_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_18_io_to_pes_5_out_bits = PE_128_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_18_io_to_pes_6_out_valid = PE_150_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_18_io_to_pes_6_out_bits = PE_150_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_18_io_to_pes_7_out_valid = PE_172_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_18_io_to_pes_7_out_bits = PE_172_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_18_io_to_pes_8_out_valid = PE_194_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_18_io_to_pes_8_out_bits = PE_194_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_18_io_to_pes_9_out_valid = PE_216_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_18_io_to_pes_9_out_bits = PE_216_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_18_io_to_pes_10_out_valid = PE_238_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_18_io_to_pes_10_out_bits = PE_238_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_18_io_to_pes_11_out_valid = PE_260_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_18_io_to_pes_11_out_bits = PE_260_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_18_io_to_pes_12_out_valid = PE_282_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_18_io_to_pes_12_out_bits = PE_282_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_18_io_to_pes_13_out_valid = PE_304_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_18_io_to_pes_13_out_bits = PE_304_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_18_io_to_pes_14_out_valid = PE_326_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_18_io_to_pes_14_out_bits = PE_326_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_18_io_to_pes_15_out_valid = PE_348_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_18_io_to_pes_15_out_bits = PE_348_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_18_io_to_pes_16_out_valid = PE_370_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_18_io_to_pes_16_out_bits = PE_370_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_18_io_to_pes_17_out_valid = PE_392_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_18_io_to_pes_17_out_bits = PE_392_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_18_io_to_pes_18_out_valid = PE_414_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_18_io_to_pes_18_out_bits = PE_414_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_18_io_to_pes_19_out_valid = PE_436_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_18_io_to_pes_19_out_bits = PE_436_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_18_io_to_pes_20_out_valid = PE_458_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_18_io_to_pes_20_out_bits = PE_458_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_18_io_to_pes_21_out_valid = PE_480_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_18_io_to_pes_21_out_bits = PE_480_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_18_io_to_pes_22_out_valid = PE_502_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_18_io_to_pes_22_out_bits = PE_502_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_18_io_to_pes_23_out_valid = PE_524_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_18_io_to_pes_23_out_bits = PE_524_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_18_io_to_pes_24_out_valid = PE_546_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_18_io_to_pes_24_out_bits = PE_546_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_18_io_to_pes_25_out_valid = PE_568_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_18_io_to_pes_25_out_bits = PE_568_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_18_io_to_pes_26_out_valid = PE_590_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_18_io_to_pes_26_out_bits = PE_590_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_18_io_to_pes_27_out_valid = PE_612_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_18_io_to_pes_27_out_bits = PE_612_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_18_io_to_pes_28_out_valid = PE_634_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_18_io_to_pes_28_out_bits = PE_634_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_18_io_to_mem_valid = MemController_18_io_rd_data_valid; // @[pe.scala 312:29]
  assign PENetwork_18_io_to_mem_bits = MemController_18_io_rd_data_bits; // @[pe.scala 312:29]
  assign PENetwork_19_io_to_pes_0_out_valid = PE_19_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_19_io_to_pes_0_out_bits = PE_19_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_19_io_to_pes_1_out_valid = PE_41_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_19_io_to_pes_1_out_bits = PE_41_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_19_io_to_pes_2_out_valid = PE_63_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_19_io_to_pes_2_out_bits = PE_63_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_19_io_to_pes_3_out_valid = PE_85_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_19_io_to_pes_3_out_bits = PE_85_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_19_io_to_pes_4_out_valid = PE_107_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_19_io_to_pes_4_out_bits = PE_107_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_19_io_to_pes_5_out_valid = PE_129_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_19_io_to_pes_5_out_bits = PE_129_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_19_io_to_pes_6_out_valid = PE_151_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_19_io_to_pes_6_out_bits = PE_151_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_19_io_to_pes_7_out_valid = PE_173_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_19_io_to_pes_7_out_bits = PE_173_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_19_io_to_pes_8_out_valid = PE_195_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_19_io_to_pes_8_out_bits = PE_195_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_19_io_to_pes_9_out_valid = PE_217_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_19_io_to_pes_9_out_bits = PE_217_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_19_io_to_pes_10_out_valid = PE_239_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_19_io_to_pes_10_out_bits = PE_239_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_19_io_to_pes_11_out_valid = PE_261_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_19_io_to_pes_11_out_bits = PE_261_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_19_io_to_pes_12_out_valid = PE_283_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_19_io_to_pes_12_out_bits = PE_283_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_19_io_to_pes_13_out_valid = PE_305_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_19_io_to_pes_13_out_bits = PE_305_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_19_io_to_pes_14_out_valid = PE_327_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_19_io_to_pes_14_out_bits = PE_327_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_19_io_to_pes_15_out_valid = PE_349_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_19_io_to_pes_15_out_bits = PE_349_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_19_io_to_pes_16_out_valid = PE_371_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_19_io_to_pes_16_out_bits = PE_371_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_19_io_to_pes_17_out_valid = PE_393_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_19_io_to_pes_17_out_bits = PE_393_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_19_io_to_pes_18_out_valid = PE_415_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_19_io_to_pes_18_out_bits = PE_415_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_19_io_to_pes_19_out_valid = PE_437_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_19_io_to_pes_19_out_bits = PE_437_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_19_io_to_pes_20_out_valid = PE_459_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_19_io_to_pes_20_out_bits = PE_459_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_19_io_to_pes_21_out_valid = PE_481_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_19_io_to_pes_21_out_bits = PE_481_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_19_io_to_pes_22_out_valid = PE_503_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_19_io_to_pes_22_out_bits = PE_503_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_19_io_to_pes_23_out_valid = PE_525_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_19_io_to_pes_23_out_bits = PE_525_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_19_io_to_pes_24_out_valid = PE_547_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_19_io_to_pes_24_out_bits = PE_547_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_19_io_to_pes_25_out_valid = PE_569_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_19_io_to_pes_25_out_bits = PE_569_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_19_io_to_pes_26_out_valid = PE_591_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_19_io_to_pes_26_out_bits = PE_591_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_19_io_to_pes_27_out_valid = PE_613_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_19_io_to_pes_27_out_bits = PE_613_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_19_io_to_pes_28_out_valid = PE_635_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_19_io_to_pes_28_out_bits = PE_635_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_19_io_to_mem_valid = MemController_19_io_rd_data_valid; // @[pe.scala 312:29]
  assign PENetwork_19_io_to_mem_bits = MemController_19_io_rd_data_bits; // @[pe.scala 312:29]
  assign PENetwork_20_io_to_pes_0_out_valid = PE_20_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_20_io_to_pes_0_out_bits = PE_20_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_20_io_to_pes_1_out_valid = PE_42_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_20_io_to_pes_1_out_bits = PE_42_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_20_io_to_pes_2_out_valid = PE_64_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_20_io_to_pes_2_out_bits = PE_64_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_20_io_to_pes_3_out_valid = PE_86_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_20_io_to_pes_3_out_bits = PE_86_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_20_io_to_pes_4_out_valid = PE_108_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_20_io_to_pes_4_out_bits = PE_108_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_20_io_to_pes_5_out_valid = PE_130_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_20_io_to_pes_5_out_bits = PE_130_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_20_io_to_pes_6_out_valid = PE_152_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_20_io_to_pes_6_out_bits = PE_152_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_20_io_to_pes_7_out_valid = PE_174_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_20_io_to_pes_7_out_bits = PE_174_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_20_io_to_pes_8_out_valid = PE_196_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_20_io_to_pes_8_out_bits = PE_196_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_20_io_to_pes_9_out_valid = PE_218_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_20_io_to_pes_9_out_bits = PE_218_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_20_io_to_pes_10_out_valid = PE_240_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_20_io_to_pes_10_out_bits = PE_240_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_20_io_to_pes_11_out_valid = PE_262_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_20_io_to_pes_11_out_bits = PE_262_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_20_io_to_pes_12_out_valid = PE_284_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_20_io_to_pes_12_out_bits = PE_284_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_20_io_to_pes_13_out_valid = PE_306_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_20_io_to_pes_13_out_bits = PE_306_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_20_io_to_pes_14_out_valid = PE_328_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_20_io_to_pes_14_out_bits = PE_328_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_20_io_to_pes_15_out_valid = PE_350_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_20_io_to_pes_15_out_bits = PE_350_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_20_io_to_pes_16_out_valid = PE_372_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_20_io_to_pes_16_out_bits = PE_372_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_20_io_to_pes_17_out_valid = PE_394_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_20_io_to_pes_17_out_bits = PE_394_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_20_io_to_pes_18_out_valid = PE_416_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_20_io_to_pes_18_out_bits = PE_416_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_20_io_to_pes_19_out_valid = PE_438_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_20_io_to_pes_19_out_bits = PE_438_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_20_io_to_pes_20_out_valid = PE_460_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_20_io_to_pes_20_out_bits = PE_460_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_20_io_to_pes_21_out_valid = PE_482_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_20_io_to_pes_21_out_bits = PE_482_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_20_io_to_pes_22_out_valid = PE_504_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_20_io_to_pes_22_out_bits = PE_504_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_20_io_to_pes_23_out_valid = PE_526_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_20_io_to_pes_23_out_bits = PE_526_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_20_io_to_pes_24_out_valid = PE_548_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_20_io_to_pes_24_out_bits = PE_548_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_20_io_to_pes_25_out_valid = PE_570_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_20_io_to_pes_25_out_bits = PE_570_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_20_io_to_pes_26_out_valid = PE_592_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_20_io_to_pes_26_out_bits = PE_592_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_20_io_to_pes_27_out_valid = PE_614_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_20_io_to_pes_27_out_bits = PE_614_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_20_io_to_pes_28_out_valid = PE_636_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_20_io_to_pes_28_out_bits = PE_636_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_20_io_to_mem_valid = MemController_20_io_rd_data_valid; // @[pe.scala 312:29]
  assign PENetwork_20_io_to_mem_bits = MemController_20_io_rd_data_bits; // @[pe.scala 312:29]
  assign PENetwork_21_io_to_pes_0_out_valid = PE_21_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_21_io_to_pes_0_out_bits = PE_21_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_21_io_to_pes_1_out_valid = PE_43_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_21_io_to_pes_1_out_bits = PE_43_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_21_io_to_pes_2_out_valid = PE_65_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_21_io_to_pes_2_out_bits = PE_65_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_21_io_to_pes_3_out_valid = PE_87_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_21_io_to_pes_3_out_bits = PE_87_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_21_io_to_pes_4_out_valid = PE_109_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_21_io_to_pes_4_out_bits = PE_109_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_21_io_to_pes_5_out_valid = PE_131_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_21_io_to_pes_5_out_bits = PE_131_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_21_io_to_pes_6_out_valid = PE_153_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_21_io_to_pes_6_out_bits = PE_153_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_21_io_to_pes_7_out_valid = PE_175_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_21_io_to_pes_7_out_bits = PE_175_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_21_io_to_pes_8_out_valid = PE_197_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_21_io_to_pes_8_out_bits = PE_197_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_21_io_to_pes_9_out_valid = PE_219_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_21_io_to_pes_9_out_bits = PE_219_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_21_io_to_pes_10_out_valid = PE_241_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_21_io_to_pes_10_out_bits = PE_241_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_21_io_to_pes_11_out_valid = PE_263_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_21_io_to_pes_11_out_bits = PE_263_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_21_io_to_pes_12_out_valid = PE_285_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_21_io_to_pes_12_out_bits = PE_285_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_21_io_to_pes_13_out_valid = PE_307_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_21_io_to_pes_13_out_bits = PE_307_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_21_io_to_pes_14_out_valid = PE_329_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_21_io_to_pes_14_out_bits = PE_329_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_21_io_to_pes_15_out_valid = PE_351_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_21_io_to_pes_15_out_bits = PE_351_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_21_io_to_pes_16_out_valid = PE_373_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_21_io_to_pes_16_out_bits = PE_373_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_21_io_to_pes_17_out_valid = PE_395_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_21_io_to_pes_17_out_bits = PE_395_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_21_io_to_pes_18_out_valid = PE_417_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_21_io_to_pes_18_out_bits = PE_417_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_21_io_to_pes_19_out_valid = PE_439_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_21_io_to_pes_19_out_bits = PE_439_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_21_io_to_pes_20_out_valid = PE_461_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_21_io_to_pes_20_out_bits = PE_461_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_21_io_to_pes_21_out_valid = PE_483_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_21_io_to_pes_21_out_bits = PE_483_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_21_io_to_pes_22_out_valid = PE_505_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_21_io_to_pes_22_out_bits = PE_505_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_21_io_to_pes_23_out_valid = PE_527_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_21_io_to_pes_23_out_bits = PE_527_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_21_io_to_pes_24_out_valid = PE_549_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_21_io_to_pes_24_out_bits = PE_549_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_21_io_to_pes_25_out_valid = PE_571_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_21_io_to_pes_25_out_bits = PE_571_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_21_io_to_pes_26_out_valid = PE_593_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_21_io_to_pes_26_out_bits = PE_593_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_21_io_to_pes_27_out_valid = PE_615_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_21_io_to_pes_27_out_bits = PE_615_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_21_io_to_pes_28_out_valid = PE_637_io_data_0_out_valid; // @[pe.scala 263:36]
  assign PENetwork_21_io_to_pes_28_out_bits = PE_637_io_data_0_out_bits; // @[pe.scala 263:36]
  assign PENetwork_21_io_to_mem_valid = MemController_21_io_rd_data_valid; // @[pe.scala 312:29]
  assign PENetwork_21_io_to_mem_bits = MemController_21_io_rd_data_bits; // @[pe.scala 312:29]
  assign PENetwork_22_io_to_pes_0_out_valid = PE_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_22_io_to_pes_0_out_bits = PE_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_22_io_to_pes_1_out_valid = PE_1_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_22_io_to_pes_1_out_bits = PE_1_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_22_io_to_pes_2_out_valid = PE_2_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_22_io_to_pes_2_out_bits = PE_2_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_22_io_to_pes_3_out_valid = PE_3_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_22_io_to_pes_3_out_bits = PE_3_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_22_io_to_pes_4_out_valid = PE_4_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_22_io_to_pes_4_out_bits = PE_4_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_22_io_to_pes_5_out_valid = PE_5_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_22_io_to_pes_5_out_bits = PE_5_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_22_io_to_pes_6_out_valid = PE_6_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_22_io_to_pes_6_out_bits = PE_6_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_22_io_to_pes_7_out_valid = PE_7_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_22_io_to_pes_7_out_bits = PE_7_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_22_io_to_pes_8_out_valid = PE_8_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_22_io_to_pes_8_out_bits = PE_8_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_22_io_to_pes_9_out_valid = PE_9_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_22_io_to_pes_9_out_bits = PE_9_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_22_io_to_pes_10_out_valid = PE_10_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_22_io_to_pes_10_out_bits = PE_10_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_22_io_to_pes_11_out_valid = PE_11_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_22_io_to_pes_11_out_bits = PE_11_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_22_io_to_pes_12_out_valid = PE_12_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_22_io_to_pes_12_out_bits = PE_12_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_22_io_to_pes_13_out_valid = PE_13_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_22_io_to_pes_13_out_bits = PE_13_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_22_io_to_pes_14_out_valid = PE_14_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_22_io_to_pes_14_out_bits = PE_14_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_22_io_to_pes_15_out_valid = PE_15_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_22_io_to_pes_15_out_bits = PE_15_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_22_io_to_pes_16_out_valid = PE_16_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_22_io_to_pes_16_out_bits = PE_16_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_22_io_to_pes_17_out_valid = PE_17_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_22_io_to_pes_17_out_bits = PE_17_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_22_io_to_pes_18_out_valid = PE_18_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_22_io_to_pes_18_out_bits = PE_18_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_22_io_to_pes_19_out_valid = PE_19_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_22_io_to_pes_19_out_bits = PE_19_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_22_io_to_pes_20_out_valid = PE_20_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_22_io_to_pes_20_out_bits = PE_20_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_22_io_to_mem_valid = MemController_22_io_rd_data_valid; // @[pe.scala 312:29]
  assign PENetwork_22_io_to_mem_bits = MemController_22_io_rd_data_bits; // @[pe.scala 312:29]
  assign PENetwork_23_io_to_pes_0_out_valid = PE_22_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_23_io_to_pes_0_out_bits = PE_22_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_23_io_to_pes_1_out_valid = PE_23_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_23_io_to_pes_1_out_bits = PE_23_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_23_io_to_pes_2_out_valid = PE_24_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_23_io_to_pes_2_out_bits = PE_24_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_23_io_to_pes_3_out_valid = PE_25_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_23_io_to_pes_3_out_bits = PE_25_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_23_io_to_pes_4_out_valid = PE_26_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_23_io_to_pes_4_out_bits = PE_26_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_23_io_to_pes_5_out_valid = PE_27_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_23_io_to_pes_5_out_bits = PE_27_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_23_io_to_pes_6_out_valid = PE_28_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_23_io_to_pes_6_out_bits = PE_28_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_23_io_to_pes_7_out_valid = PE_29_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_23_io_to_pes_7_out_bits = PE_29_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_23_io_to_pes_8_out_valid = PE_30_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_23_io_to_pes_8_out_bits = PE_30_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_23_io_to_pes_9_out_valid = PE_31_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_23_io_to_pes_9_out_bits = PE_31_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_23_io_to_pes_10_out_valid = PE_32_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_23_io_to_pes_10_out_bits = PE_32_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_23_io_to_pes_11_out_valid = PE_33_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_23_io_to_pes_11_out_bits = PE_33_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_23_io_to_pes_12_out_valid = PE_34_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_23_io_to_pes_12_out_bits = PE_34_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_23_io_to_pes_13_out_valid = PE_35_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_23_io_to_pes_13_out_bits = PE_35_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_23_io_to_pes_14_out_valid = PE_36_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_23_io_to_pes_14_out_bits = PE_36_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_23_io_to_pes_15_out_valid = PE_37_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_23_io_to_pes_15_out_bits = PE_37_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_23_io_to_pes_16_out_valid = PE_38_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_23_io_to_pes_16_out_bits = PE_38_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_23_io_to_pes_17_out_valid = PE_39_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_23_io_to_pes_17_out_bits = PE_39_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_23_io_to_pes_18_out_valid = PE_40_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_23_io_to_pes_18_out_bits = PE_40_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_23_io_to_pes_19_out_valid = PE_41_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_23_io_to_pes_19_out_bits = PE_41_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_23_io_to_pes_20_out_valid = PE_42_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_23_io_to_pes_20_out_bits = PE_42_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_23_io_to_mem_valid = MemController_23_io_rd_data_valid; // @[pe.scala 312:29]
  assign PENetwork_23_io_to_mem_bits = MemController_23_io_rd_data_bits; // @[pe.scala 312:29]
  assign PENetwork_24_io_to_pes_0_out_valid = PE_44_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_24_io_to_pes_0_out_bits = PE_44_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_24_io_to_pes_1_out_valid = PE_45_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_24_io_to_pes_1_out_bits = PE_45_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_24_io_to_pes_2_out_valid = PE_46_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_24_io_to_pes_2_out_bits = PE_46_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_24_io_to_pes_3_out_valid = PE_47_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_24_io_to_pes_3_out_bits = PE_47_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_24_io_to_pes_4_out_valid = PE_48_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_24_io_to_pes_4_out_bits = PE_48_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_24_io_to_pes_5_out_valid = PE_49_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_24_io_to_pes_5_out_bits = PE_49_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_24_io_to_pes_6_out_valid = PE_50_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_24_io_to_pes_6_out_bits = PE_50_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_24_io_to_pes_7_out_valid = PE_51_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_24_io_to_pes_7_out_bits = PE_51_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_24_io_to_pes_8_out_valid = PE_52_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_24_io_to_pes_8_out_bits = PE_52_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_24_io_to_pes_9_out_valid = PE_53_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_24_io_to_pes_9_out_bits = PE_53_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_24_io_to_pes_10_out_valid = PE_54_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_24_io_to_pes_10_out_bits = PE_54_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_24_io_to_pes_11_out_valid = PE_55_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_24_io_to_pes_11_out_bits = PE_55_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_24_io_to_pes_12_out_valid = PE_56_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_24_io_to_pes_12_out_bits = PE_56_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_24_io_to_pes_13_out_valid = PE_57_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_24_io_to_pes_13_out_bits = PE_57_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_24_io_to_pes_14_out_valid = PE_58_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_24_io_to_pes_14_out_bits = PE_58_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_24_io_to_pes_15_out_valid = PE_59_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_24_io_to_pes_15_out_bits = PE_59_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_24_io_to_pes_16_out_valid = PE_60_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_24_io_to_pes_16_out_bits = PE_60_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_24_io_to_pes_17_out_valid = PE_61_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_24_io_to_pes_17_out_bits = PE_61_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_24_io_to_pes_18_out_valid = PE_62_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_24_io_to_pes_18_out_bits = PE_62_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_24_io_to_pes_19_out_valid = PE_63_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_24_io_to_pes_19_out_bits = PE_63_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_24_io_to_pes_20_out_valid = PE_64_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_24_io_to_pes_20_out_bits = PE_64_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_24_io_to_mem_valid = MemController_24_io_rd_data_valid; // @[pe.scala 312:29]
  assign PENetwork_24_io_to_mem_bits = MemController_24_io_rd_data_bits; // @[pe.scala 312:29]
  assign PENetwork_25_io_to_pes_0_out_valid = PE_66_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_25_io_to_pes_0_out_bits = PE_66_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_25_io_to_pes_1_out_valid = PE_67_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_25_io_to_pes_1_out_bits = PE_67_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_25_io_to_pes_2_out_valid = PE_68_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_25_io_to_pes_2_out_bits = PE_68_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_25_io_to_pes_3_out_valid = PE_69_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_25_io_to_pes_3_out_bits = PE_69_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_25_io_to_pes_4_out_valid = PE_70_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_25_io_to_pes_4_out_bits = PE_70_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_25_io_to_pes_5_out_valid = PE_71_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_25_io_to_pes_5_out_bits = PE_71_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_25_io_to_pes_6_out_valid = PE_72_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_25_io_to_pes_6_out_bits = PE_72_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_25_io_to_pes_7_out_valid = PE_73_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_25_io_to_pes_7_out_bits = PE_73_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_25_io_to_pes_8_out_valid = PE_74_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_25_io_to_pes_8_out_bits = PE_74_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_25_io_to_pes_9_out_valid = PE_75_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_25_io_to_pes_9_out_bits = PE_75_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_25_io_to_pes_10_out_valid = PE_76_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_25_io_to_pes_10_out_bits = PE_76_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_25_io_to_pes_11_out_valid = PE_77_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_25_io_to_pes_11_out_bits = PE_77_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_25_io_to_pes_12_out_valid = PE_78_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_25_io_to_pes_12_out_bits = PE_78_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_25_io_to_pes_13_out_valid = PE_79_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_25_io_to_pes_13_out_bits = PE_79_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_25_io_to_pes_14_out_valid = PE_80_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_25_io_to_pes_14_out_bits = PE_80_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_25_io_to_pes_15_out_valid = PE_81_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_25_io_to_pes_15_out_bits = PE_81_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_25_io_to_pes_16_out_valid = PE_82_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_25_io_to_pes_16_out_bits = PE_82_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_25_io_to_pes_17_out_valid = PE_83_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_25_io_to_pes_17_out_bits = PE_83_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_25_io_to_pes_18_out_valid = PE_84_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_25_io_to_pes_18_out_bits = PE_84_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_25_io_to_pes_19_out_valid = PE_85_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_25_io_to_pes_19_out_bits = PE_85_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_25_io_to_pes_20_out_valid = PE_86_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_25_io_to_pes_20_out_bits = PE_86_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_25_io_to_mem_valid = MemController_25_io_rd_data_valid; // @[pe.scala 312:29]
  assign PENetwork_25_io_to_mem_bits = MemController_25_io_rd_data_bits; // @[pe.scala 312:29]
  assign PENetwork_26_io_to_pes_0_out_valid = PE_88_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_26_io_to_pes_0_out_bits = PE_88_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_26_io_to_pes_1_out_valid = PE_89_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_26_io_to_pes_1_out_bits = PE_89_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_26_io_to_pes_2_out_valid = PE_90_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_26_io_to_pes_2_out_bits = PE_90_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_26_io_to_pes_3_out_valid = PE_91_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_26_io_to_pes_3_out_bits = PE_91_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_26_io_to_pes_4_out_valid = PE_92_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_26_io_to_pes_4_out_bits = PE_92_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_26_io_to_pes_5_out_valid = PE_93_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_26_io_to_pes_5_out_bits = PE_93_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_26_io_to_pes_6_out_valid = PE_94_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_26_io_to_pes_6_out_bits = PE_94_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_26_io_to_pes_7_out_valid = PE_95_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_26_io_to_pes_7_out_bits = PE_95_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_26_io_to_pes_8_out_valid = PE_96_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_26_io_to_pes_8_out_bits = PE_96_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_26_io_to_pes_9_out_valid = PE_97_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_26_io_to_pes_9_out_bits = PE_97_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_26_io_to_pes_10_out_valid = PE_98_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_26_io_to_pes_10_out_bits = PE_98_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_26_io_to_pes_11_out_valid = PE_99_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_26_io_to_pes_11_out_bits = PE_99_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_26_io_to_pes_12_out_valid = PE_100_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_26_io_to_pes_12_out_bits = PE_100_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_26_io_to_pes_13_out_valid = PE_101_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_26_io_to_pes_13_out_bits = PE_101_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_26_io_to_pes_14_out_valid = PE_102_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_26_io_to_pes_14_out_bits = PE_102_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_26_io_to_pes_15_out_valid = PE_103_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_26_io_to_pes_15_out_bits = PE_103_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_26_io_to_pes_16_out_valid = PE_104_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_26_io_to_pes_16_out_bits = PE_104_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_26_io_to_pes_17_out_valid = PE_105_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_26_io_to_pes_17_out_bits = PE_105_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_26_io_to_pes_18_out_valid = PE_106_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_26_io_to_pes_18_out_bits = PE_106_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_26_io_to_pes_19_out_valid = PE_107_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_26_io_to_pes_19_out_bits = PE_107_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_26_io_to_pes_20_out_valid = PE_108_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_26_io_to_pes_20_out_bits = PE_108_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_26_io_to_mem_valid = MemController_26_io_rd_data_valid; // @[pe.scala 312:29]
  assign PENetwork_26_io_to_mem_bits = MemController_26_io_rd_data_bits; // @[pe.scala 312:29]
  assign PENetwork_27_io_to_pes_0_out_valid = PE_110_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_27_io_to_pes_0_out_bits = PE_110_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_27_io_to_pes_1_out_valid = PE_111_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_27_io_to_pes_1_out_bits = PE_111_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_27_io_to_pes_2_out_valid = PE_112_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_27_io_to_pes_2_out_bits = PE_112_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_27_io_to_pes_3_out_valid = PE_113_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_27_io_to_pes_3_out_bits = PE_113_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_27_io_to_pes_4_out_valid = PE_114_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_27_io_to_pes_4_out_bits = PE_114_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_27_io_to_pes_5_out_valid = PE_115_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_27_io_to_pes_5_out_bits = PE_115_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_27_io_to_pes_6_out_valid = PE_116_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_27_io_to_pes_6_out_bits = PE_116_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_27_io_to_pes_7_out_valid = PE_117_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_27_io_to_pes_7_out_bits = PE_117_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_27_io_to_pes_8_out_valid = PE_118_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_27_io_to_pes_8_out_bits = PE_118_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_27_io_to_pes_9_out_valid = PE_119_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_27_io_to_pes_9_out_bits = PE_119_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_27_io_to_pes_10_out_valid = PE_120_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_27_io_to_pes_10_out_bits = PE_120_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_27_io_to_pes_11_out_valid = PE_121_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_27_io_to_pes_11_out_bits = PE_121_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_27_io_to_pes_12_out_valid = PE_122_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_27_io_to_pes_12_out_bits = PE_122_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_27_io_to_pes_13_out_valid = PE_123_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_27_io_to_pes_13_out_bits = PE_123_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_27_io_to_pes_14_out_valid = PE_124_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_27_io_to_pes_14_out_bits = PE_124_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_27_io_to_pes_15_out_valid = PE_125_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_27_io_to_pes_15_out_bits = PE_125_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_27_io_to_pes_16_out_valid = PE_126_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_27_io_to_pes_16_out_bits = PE_126_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_27_io_to_pes_17_out_valid = PE_127_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_27_io_to_pes_17_out_bits = PE_127_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_27_io_to_pes_18_out_valid = PE_128_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_27_io_to_pes_18_out_bits = PE_128_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_27_io_to_pes_19_out_valid = PE_129_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_27_io_to_pes_19_out_bits = PE_129_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_27_io_to_pes_20_out_valid = PE_130_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_27_io_to_pes_20_out_bits = PE_130_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_27_io_to_mem_valid = MemController_27_io_rd_data_valid; // @[pe.scala 312:29]
  assign PENetwork_27_io_to_mem_bits = MemController_27_io_rd_data_bits; // @[pe.scala 312:29]
  assign PENetwork_28_io_to_pes_0_out_valid = PE_132_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_28_io_to_pes_0_out_bits = PE_132_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_28_io_to_pes_1_out_valid = PE_133_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_28_io_to_pes_1_out_bits = PE_133_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_28_io_to_pes_2_out_valid = PE_134_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_28_io_to_pes_2_out_bits = PE_134_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_28_io_to_pes_3_out_valid = PE_135_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_28_io_to_pes_3_out_bits = PE_135_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_28_io_to_pes_4_out_valid = PE_136_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_28_io_to_pes_4_out_bits = PE_136_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_28_io_to_pes_5_out_valid = PE_137_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_28_io_to_pes_5_out_bits = PE_137_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_28_io_to_pes_6_out_valid = PE_138_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_28_io_to_pes_6_out_bits = PE_138_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_28_io_to_pes_7_out_valid = PE_139_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_28_io_to_pes_7_out_bits = PE_139_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_28_io_to_pes_8_out_valid = PE_140_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_28_io_to_pes_8_out_bits = PE_140_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_28_io_to_pes_9_out_valid = PE_141_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_28_io_to_pes_9_out_bits = PE_141_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_28_io_to_pes_10_out_valid = PE_142_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_28_io_to_pes_10_out_bits = PE_142_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_28_io_to_pes_11_out_valid = PE_143_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_28_io_to_pes_11_out_bits = PE_143_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_28_io_to_pes_12_out_valid = PE_144_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_28_io_to_pes_12_out_bits = PE_144_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_28_io_to_pes_13_out_valid = PE_145_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_28_io_to_pes_13_out_bits = PE_145_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_28_io_to_pes_14_out_valid = PE_146_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_28_io_to_pes_14_out_bits = PE_146_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_28_io_to_pes_15_out_valid = PE_147_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_28_io_to_pes_15_out_bits = PE_147_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_28_io_to_pes_16_out_valid = PE_148_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_28_io_to_pes_16_out_bits = PE_148_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_28_io_to_pes_17_out_valid = PE_149_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_28_io_to_pes_17_out_bits = PE_149_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_28_io_to_pes_18_out_valid = PE_150_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_28_io_to_pes_18_out_bits = PE_150_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_28_io_to_pes_19_out_valid = PE_151_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_28_io_to_pes_19_out_bits = PE_151_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_28_io_to_pes_20_out_valid = PE_152_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_28_io_to_pes_20_out_bits = PE_152_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_28_io_to_mem_valid = MemController_28_io_rd_data_valid; // @[pe.scala 312:29]
  assign PENetwork_28_io_to_mem_bits = MemController_28_io_rd_data_bits; // @[pe.scala 312:29]
  assign PENetwork_29_io_to_pes_0_out_valid = PE_154_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_29_io_to_pes_0_out_bits = PE_154_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_29_io_to_pes_1_out_valid = PE_155_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_29_io_to_pes_1_out_bits = PE_155_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_29_io_to_pes_2_out_valid = PE_156_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_29_io_to_pes_2_out_bits = PE_156_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_29_io_to_pes_3_out_valid = PE_157_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_29_io_to_pes_3_out_bits = PE_157_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_29_io_to_pes_4_out_valid = PE_158_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_29_io_to_pes_4_out_bits = PE_158_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_29_io_to_pes_5_out_valid = PE_159_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_29_io_to_pes_5_out_bits = PE_159_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_29_io_to_pes_6_out_valid = PE_160_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_29_io_to_pes_6_out_bits = PE_160_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_29_io_to_pes_7_out_valid = PE_161_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_29_io_to_pes_7_out_bits = PE_161_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_29_io_to_pes_8_out_valid = PE_162_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_29_io_to_pes_8_out_bits = PE_162_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_29_io_to_pes_9_out_valid = PE_163_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_29_io_to_pes_9_out_bits = PE_163_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_29_io_to_pes_10_out_valid = PE_164_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_29_io_to_pes_10_out_bits = PE_164_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_29_io_to_pes_11_out_valid = PE_165_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_29_io_to_pes_11_out_bits = PE_165_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_29_io_to_pes_12_out_valid = PE_166_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_29_io_to_pes_12_out_bits = PE_166_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_29_io_to_pes_13_out_valid = PE_167_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_29_io_to_pes_13_out_bits = PE_167_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_29_io_to_pes_14_out_valid = PE_168_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_29_io_to_pes_14_out_bits = PE_168_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_29_io_to_pes_15_out_valid = PE_169_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_29_io_to_pes_15_out_bits = PE_169_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_29_io_to_pes_16_out_valid = PE_170_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_29_io_to_pes_16_out_bits = PE_170_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_29_io_to_pes_17_out_valid = PE_171_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_29_io_to_pes_17_out_bits = PE_171_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_29_io_to_pes_18_out_valid = PE_172_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_29_io_to_pes_18_out_bits = PE_172_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_29_io_to_pes_19_out_valid = PE_173_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_29_io_to_pes_19_out_bits = PE_173_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_29_io_to_pes_20_out_valid = PE_174_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_29_io_to_pes_20_out_bits = PE_174_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_29_io_to_mem_valid = MemController_29_io_rd_data_valid; // @[pe.scala 312:29]
  assign PENetwork_29_io_to_mem_bits = MemController_29_io_rd_data_bits; // @[pe.scala 312:29]
  assign PENetwork_30_io_to_pes_0_out_valid = PE_176_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_30_io_to_pes_0_out_bits = PE_176_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_30_io_to_pes_1_out_valid = PE_177_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_30_io_to_pes_1_out_bits = PE_177_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_30_io_to_pes_2_out_valid = PE_178_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_30_io_to_pes_2_out_bits = PE_178_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_30_io_to_pes_3_out_valid = PE_179_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_30_io_to_pes_3_out_bits = PE_179_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_30_io_to_pes_4_out_valid = PE_180_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_30_io_to_pes_4_out_bits = PE_180_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_30_io_to_pes_5_out_valid = PE_181_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_30_io_to_pes_5_out_bits = PE_181_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_30_io_to_pes_6_out_valid = PE_182_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_30_io_to_pes_6_out_bits = PE_182_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_30_io_to_pes_7_out_valid = PE_183_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_30_io_to_pes_7_out_bits = PE_183_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_30_io_to_pes_8_out_valid = PE_184_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_30_io_to_pes_8_out_bits = PE_184_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_30_io_to_pes_9_out_valid = PE_185_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_30_io_to_pes_9_out_bits = PE_185_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_30_io_to_pes_10_out_valid = PE_186_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_30_io_to_pes_10_out_bits = PE_186_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_30_io_to_pes_11_out_valid = PE_187_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_30_io_to_pes_11_out_bits = PE_187_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_30_io_to_pes_12_out_valid = PE_188_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_30_io_to_pes_12_out_bits = PE_188_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_30_io_to_pes_13_out_valid = PE_189_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_30_io_to_pes_13_out_bits = PE_189_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_30_io_to_pes_14_out_valid = PE_190_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_30_io_to_pes_14_out_bits = PE_190_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_30_io_to_pes_15_out_valid = PE_191_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_30_io_to_pes_15_out_bits = PE_191_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_30_io_to_pes_16_out_valid = PE_192_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_30_io_to_pes_16_out_bits = PE_192_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_30_io_to_pes_17_out_valid = PE_193_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_30_io_to_pes_17_out_bits = PE_193_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_30_io_to_pes_18_out_valid = PE_194_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_30_io_to_pes_18_out_bits = PE_194_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_30_io_to_pes_19_out_valid = PE_195_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_30_io_to_pes_19_out_bits = PE_195_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_30_io_to_pes_20_out_valid = PE_196_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_30_io_to_pes_20_out_bits = PE_196_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_30_io_to_mem_valid = MemController_30_io_rd_data_valid; // @[pe.scala 312:29]
  assign PENetwork_30_io_to_mem_bits = MemController_30_io_rd_data_bits; // @[pe.scala 312:29]
  assign PENetwork_31_io_to_pes_0_out_valid = PE_198_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_31_io_to_pes_0_out_bits = PE_198_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_31_io_to_pes_1_out_valid = PE_199_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_31_io_to_pes_1_out_bits = PE_199_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_31_io_to_pes_2_out_valid = PE_200_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_31_io_to_pes_2_out_bits = PE_200_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_31_io_to_pes_3_out_valid = PE_201_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_31_io_to_pes_3_out_bits = PE_201_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_31_io_to_pes_4_out_valid = PE_202_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_31_io_to_pes_4_out_bits = PE_202_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_31_io_to_pes_5_out_valid = PE_203_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_31_io_to_pes_5_out_bits = PE_203_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_31_io_to_pes_6_out_valid = PE_204_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_31_io_to_pes_6_out_bits = PE_204_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_31_io_to_pes_7_out_valid = PE_205_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_31_io_to_pes_7_out_bits = PE_205_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_31_io_to_pes_8_out_valid = PE_206_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_31_io_to_pes_8_out_bits = PE_206_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_31_io_to_pes_9_out_valid = PE_207_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_31_io_to_pes_9_out_bits = PE_207_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_31_io_to_pes_10_out_valid = PE_208_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_31_io_to_pes_10_out_bits = PE_208_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_31_io_to_pes_11_out_valid = PE_209_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_31_io_to_pes_11_out_bits = PE_209_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_31_io_to_pes_12_out_valid = PE_210_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_31_io_to_pes_12_out_bits = PE_210_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_31_io_to_pes_13_out_valid = PE_211_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_31_io_to_pes_13_out_bits = PE_211_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_31_io_to_pes_14_out_valid = PE_212_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_31_io_to_pes_14_out_bits = PE_212_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_31_io_to_pes_15_out_valid = PE_213_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_31_io_to_pes_15_out_bits = PE_213_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_31_io_to_pes_16_out_valid = PE_214_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_31_io_to_pes_16_out_bits = PE_214_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_31_io_to_pes_17_out_valid = PE_215_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_31_io_to_pes_17_out_bits = PE_215_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_31_io_to_pes_18_out_valid = PE_216_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_31_io_to_pes_18_out_bits = PE_216_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_31_io_to_pes_19_out_valid = PE_217_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_31_io_to_pes_19_out_bits = PE_217_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_31_io_to_pes_20_out_valid = PE_218_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_31_io_to_pes_20_out_bits = PE_218_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_31_io_to_mem_valid = MemController_31_io_rd_data_valid; // @[pe.scala 312:29]
  assign PENetwork_31_io_to_mem_bits = MemController_31_io_rd_data_bits; // @[pe.scala 312:29]
  assign PENetwork_32_io_to_pes_0_out_valid = PE_220_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_32_io_to_pes_0_out_bits = PE_220_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_32_io_to_pes_1_out_valid = PE_221_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_32_io_to_pes_1_out_bits = PE_221_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_32_io_to_pes_2_out_valid = PE_222_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_32_io_to_pes_2_out_bits = PE_222_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_32_io_to_pes_3_out_valid = PE_223_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_32_io_to_pes_3_out_bits = PE_223_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_32_io_to_pes_4_out_valid = PE_224_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_32_io_to_pes_4_out_bits = PE_224_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_32_io_to_pes_5_out_valid = PE_225_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_32_io_to_pes_5_out_bits = PE_225_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_32_io_to_pes_6_out_valid = PE_226_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_32_io_to_pes_6_out_bits = PE_226_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_32_io_to_pes_7_out_valid = PE_227_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_32_io_to_pes_7_out_bits = PE_227_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_32_io_to_pes_8_out_valid = PE_228_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_32_io_to_pes_8_out_bits = PE_228_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_32_io_to_pes_9_out_valid = PE_229_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_32_io_to_pes_9_out_bits = PE_229_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_32_io_to_pes_10_out_valid = PE_230_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_32_io_to_pes_10_out_bits = PE_230_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_32_io_to_pes_11_out_valid = PE_231_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_32_io_to_pes_11_out_bits = PE_231_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_32_io_to_pes_12_out_valid = PE_232_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_32_io_to_pes_12_out_bits = PE_232_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_32_io_to_pes_13_out_valid = PE_233_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_32_io_to_pes_13_out_bits = PE_233_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_32_io_to_pes_14_out_valid = PE_234_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_32_io_to_pes_14_out_bits = PE_234_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_32_io_to_pes_15_out_valid = PE_235_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_32_io_to_pes_15_out_bits = PE_235_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_32_io_to_pes_16_out_valid = PE_236_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_32_io_to_pes_16_out_bits = PE_236_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_32_io_to_pes_17_out_valid = PE_237_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_32_io_to_pes_17_out_bits = PE_237_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_32_io_to_pes_18_out_valid = PE_238_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_32_io_to_pes_18_out_bits = PE_238_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_32_io_to_pes_19_out_valid = PE_239_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_32_io_to_pes_19_out_bits = PE_239_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_32_io_to_pes_20_out_valid = PE_240_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_32_io_to_pes_20_out_bits = PE_240_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_32_io_to_mem_valid = MemController_32_io_rd_data_valid; // @[pe.scala 312:29]
  assign PENetwork_32_io_to_mem_bits = MemController_32_io_rd_data_bits; // @[pe.scala 312:29]
  assign PENetwork_33_io_to_pes_0_out_valid = PE_242_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_33_io_to_pes_0_out_bits = PE_242_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_33_io_to_pes_1_out_valid = PE_243_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_33_io_to_pes_1_out_bits = PE_243_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_33_io_to_pes_2_out_valid = PE_244_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_33_io_to_pes_2_out_bits = PE_244_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_33_io_to_pes_3_out_valid = PE_245_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_33_io_to_pes_3_out_bits = PE_245_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_33_io_to_pes_4_out_valid = PE_246_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_33_io_to_pes_4_out_bits = PE_246_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_33_io_to_pes_5_out_valid = PE_247_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_33_io_to_pes_5_out_bits = PE_247_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_33_io_to_pes_6_out_valid = PE_248_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_33_io_to_pes_6_out_bits = PE_248_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_33_io_to_pes_7_out_valid = PE_249_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_33_io_to_pes_7_out_bits = PE_249_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_33_io_to_pes_8_out_valid = PE_250_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_33_io_to_pes_8_out_bits = PE_250_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_33_io_to_pes_9_out_valid = PE_251_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_33_io_to_pes_9_out_bits = PE_251_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_33_io_to_pes_10_out_valid = PE_252_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_33_io_to_pes_10_out_bits = PE_252_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_33_io_to_pes_11_out_valid = PE_253_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_33_io_to_pes_11_out_bits = PE_253_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_33_io_to_pes_12_out_valid = PE_254_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_33_io_to_pes_12_out_bits = PE_254_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_33_io_to_pes_13_out_valid = PE_255_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_33_io_to_pes_13_out_bits = PE_255_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_33_io_to_pes_14_out_valid = PE_256_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_33_io_to_pes_14_out_bits = PE_256_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_33_io_to_pes_15_out_valid = PE_257_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_33_io_to_pes_15_out_bits = PE_257_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_33_io_to_pes_16_out_valid = PE_258_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_33_io_to_pes_16_out_bits = PE_258_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_33_io_to_pes_17_out_valid = PE_259_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_33_io_to_pes_17_out_bits = PE_259_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_33_io_to_pes_18_out_valid = PE_260_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_33_io_to_pes_18_out_bits = PE_260_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_33_io_to_pes_19_out_valid = PE_261_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_33_io_to_pes_19_out_bits = PE_261_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_33_io_to_pes_20_out_valid = PE_262_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_33_io_to_pes_20_out_bits = PE_262_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_33_io_to_mem_valid = MemController_33_io_rd_data_valid; // @[pe.scala 312:29]
  assign PENetwork_33_io_to_mem_bits = MemController_33_io_rd_data_bits; // @[pe.scala 312:29]
  assign PENetwork_34_io_to_pes_0_out_valid = PE_264_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_34_io_to_pes_0_out_bits = PE_264_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_34_io_to_pes_1_out_valid = PE_265_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_34_io_to_pes_1_out_bits = PE_265_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_34_io_to_pes_2_out_valid = PE_266_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_34_io_to_pes_2_out_bits = PE_266_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_34_io_to_pes_3_out_valid = PE_267_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_34_io_to_pes_3_out_bits = PE_267_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_34_io_to_pes_4_out_valid = PE_268_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_34_io_to_pes_4_out_bits = PE_268_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_34_io_to_pes_5_out_valid = PE_269_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_34_io_to_pes_5_out_bits = PE_269_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_34_io_to_pes_6_out_valid = PE_270_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_34_io_to_pes_6_out_bits = PE_270_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_34_io_to_pes_7_out_valid = PE_271_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_34_io_to_pes_7_out_bits = PE_271_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_34_io_to_pes_8_out_valid = PE_272_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_34_io_to_pes_8_out_bits = PE_272_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_34_io_to_pes_9_out_valid = PE_273_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_34_io_to_pes_9_out_bits = PE_273_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_34_io_to_pes_10_out_valid = PE_274_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_34_io_to_pes_10_out_bits = PE_274_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_34_io_to_pes_11_out_valid = PE_275_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_34_io_to_pes_11_out_bits = PE_275_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_34_io_to_pes_12_out_valid = PE_276_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_34_io_to_pes_12_out_bits = PE_276_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_34_io_to_pes_13_out_valid = PE_277_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_34_io_to_pes_13_out_bits = PE_277_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_34_io_to_pes_14_out_valid = PE_278_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_34_io_to_pes_14_out_bits = PE_278_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_34_io_to_pes_15_out_valid = PE_279_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_34_io_to_pes_15_out_bits = PE_279_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_34_io_to_pes_16_out_valid = PE_280_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_34_io_to_pes_16_out_bits = PE_280_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_34_io_to_pes_17_out_valid = PE_281_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_34_io_to_pes_17_out_bits = PE_281_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_34_io_to_pes_18_out_valid = PE_282_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_34_io_to_pes_18_out_bits = PE_282_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_34_io_to_pes_19_out_valid = PE_283_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_34_io_to_pes_19_out_bits = PE_283_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_34_io_to_pes_20_out_valid = PE_284_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_34_io_to_pes_20_out_bits = PE_284_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_34_io_to_mem_valid = MemController_34_io_rd_data_valid; // @[pe.scala 312:29]
  assign PENetwork_34_io_to_mem_bits = MemController_34_io_rd_data_bits; // @[pe.scala 312:29]
  assign PENetwork_35_io_to_pes_0_out_valid = PE_286_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_35_io_to_pes_0_out_bits = PE_286_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_35_io_to_pes_1_out_valid = PE_287_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_35_io_to_pes_1_out_bits = PE_287_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_35_io_to_pes_2_out_valid = PE_288_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_35_io_to_pes_2_out_bits = PE_288_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_35_io_to_pes_3_out_valid = PE_289_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_35_io_to_pes_3_out_bits = PE_289_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_35_io_to_pes_4_out_valid = PE_290_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_35_io_to_pes_4_out_bits = PE_290_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_35_io_to_pes_5_out_valid = PE_291_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_35_io_to_pes_5_out_bits = PE_291_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_35_io_to_pes_6_out_valid = PE_292_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_35_io_to_pes_6_out_bits = PE_292_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_35_io_to_pes_7_out_valid = PE_293_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_35_io_to_pes_7_out_bits = PE_293_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_35_io_to_pes_8_out_valid = PE_294_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_35_io_to_pes_8_out_bits = PE_294_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_35_io_to_pes_9_out_valid = PE_295_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_35_io_to_pes_9_out_bits = PE_295_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_35_io_to_pes_10_out_valid = PE_296_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_35_io_to_pes_10_out_bits = PE_296_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_35_io_to_pes_11_out_valid = PE_297_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_35_io_to_pes_11_out_bits = PE_297_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_35_io_to_pes_12_out_valid = PE_298_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_35_io_to_pes_12_out_bits = PE_298_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_35_io_to_pes_13_out_valid = PE_299_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_35_io_to_pes_13_out_bits = PE_299_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_35_io_to_pes_14_out_valid = PE_300_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_35_io_to_pes_14_out_bits = PE_300_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_35_io_to_pes_15_out_valid = PE_301_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_35_io_to_pes_15_out_bits = PE_301_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_35_io_to_pes_16_out_valid = PE_302_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_35_io_to_pes_16_out_bits = PE_302_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_35_io_to_pes_17_out_valid = PE_303_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_35_io_to_pes_17_out_bits = PE_303_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_35_io_to_pes_18_out_valid = PE_304_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_35_io_to_pes_18_out_bits = PE_304_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_35_io_to_pes_19_out_valid = PE_305_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_35_io_to_pes_19_out_bits = PE_305_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_35_io_to_pes_20_out_valid = PE_306_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_35_io_to_pes_20_out_bits = PE_306_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_35_io_to_mem_valid = MemController_35_io_rd_data_valid; // @[pe.scala 312:29]
  assign PENetwork_35_io_to_mem_bits = MemController_35_io_rd_data_bits; // @[pe.scala 312:29]
  assign PENetwork_36_io_to_pes_0_out_valid = PE_308_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_36_io_to_pes_0_out_bits = PE_308_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_36_io_to_pes_1_out_valid = PE_309_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_36_io_to_pes_1_out_bits = PE_309_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_36_io_to_pes_2_out_valid = PE_310_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_36_io_to_pes_2_out_bits = PE_310_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_36_io_to_pes_3_out_valid = PE_311_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_36_io_to_pes_3_out_bits = PE_311_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_36_io_to_pes_4_out_valid = PE_312_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_36_io_to_pes_4_out_bits = PE_312_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_36_io_to_pes_5_out_valid = PE_313_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_36_io_to_pes_5_out_bits = PE_313_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_36_io_to_pes_6_out_valid = PE_314_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_36_io_to_pes_6_out_bits = PE_314_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_36_io_to_pes_7_out_valid = PE_315_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_36_io_to_pes_7_out_bits = PE_315_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_36_io_to_pes_8_out_valid = PE_316_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_36_io_to_pes_8_out_bits = PE_316_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_36_io_to_pes_9_out_valid = PE_317_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_36_io_to_pes_9_out_bits = PE_317_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_36_io_to_pes_10_out_valid = PE_318_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_36_io_to_pes_10_out_bits = PE_318_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_36_io_to_pes_11_out_valid = PE_319_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_36_io_to_pes_11_out_bits = PE_319_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_36_io_to_pes_12_out_valid = PE_320_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_36_io_to_pes_12_out_bits = PE_320_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_36_io_to_pes_13_out_valid = PE_321_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_36_io_to_pes_13_out_bits = PE_321_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_36_io_to_pes_14_out_valid = PE_322_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_36_io_to_pes_14_out_bits = PE_322_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_36_io_to_pes_15_out_valid = PE_323_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_36_io_to_pes_15_out_bits = PE_323_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_36_io_to_pes_16_out_valid = PE_324_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_36_io_to_pes_16_out_bits = PE_324_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_36_io_to_pes_17_out_valid = PE_325_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_36_io_to_pes_17_out_bits = PE_325_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_36_io_to_pes_18_out_valid = PE_326_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_36_io_to_pes_18_out_bits = PE_326_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_36_io_to_pes_19_out_valid = PE_327_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_36_io_to_pes_19_out_bits = PE_327_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_36_io_to_pes_20_out_valid = PE_328_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_36_io_to_pes_20_out_bits = PE_328_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_36_io_to_mem_valid = MemController_36_io_rd_data_valid; // @[pe.scala 312:29]
  assign PENetwork_36_io_to_mem_bits = MemController_36_io_rd_data_bits; // @[pe.scala 312:29]
  assign PENetwork_37_io_to_pes_0_out_valid = PE_330_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_37_io_to_pes_0_out_bits = PE_330_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_37_io_to_pes_1_out_valid = PE_331_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_37_io_to_pes_1_out_bits = PE_331_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_37_io_to_pes_2_out_valid = PE_332_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_37_io_to_pes_2_out_bits = PE_332_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_37_io_to_pes_3_out_valid = PE_333_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_37_io_to_pes_3_out_bits = PE_333_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_37_io_to_pes_4_out_valid = PE_334_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_37_io_to_pes_4_out_bits = PE_334_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_37_io_to_pes_5_out_valid = PE_335_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_37_io_to_pes_5_out_bits = PE_335_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_37_io_to_pes_6_out_valid = PE_336_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_37_io_to_pes_6_out_bits = PE_336_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_37_io_to_pes_7_out_valid = PE_337_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_37_io_to_pes_7_out_bits = PE_337_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_37_io_to_pes_8_out_valid = PE_338_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_37_io_to_pes_8_out_bits = PE_338_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_37_io_to_pes_9_out_valid = PE_339_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_37_io_to_pes_9_out_bits = PE_339_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_37_io_to_pes_10_out_valid = PE_340_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_37_io_to_pes_10_out_bits = PE_340_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_37_io_to_pes_11_out_valid = PE_341_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_37_io_to_pes_11_out_bits = PE_341_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_37_io_to_pes_12_out_valid = PE_342_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_37_io_to_pes_12_out_bits = PE_342_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_37_io_to_pes_13_out_valid = PE_343_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_37_io_to_pes_13_out_bits = PE_343_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_37_io_to_pes_14_out_valid = PE_344_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_37_io_to_pes_14_out_bits = PE_344_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_37_io_to_pes_15_out_valid = PE_345_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_37_io_to_pes_15_out_bits = PE_345_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_37_io_to_pes_16_out_valid = PE_346_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_37_io_to_pes_16_out_bits = PE_346_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_37_io_to_pes_17_out_valid = PE_347_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_37_io_to_pes_17_out_bits = PE_347_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_37_io_to_pes_18_out_valid = PE_348_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_37_io_to_pes_18_out_bits = PE_348_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_37_io_to_pes_19_out_valid = PE_349_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_37_io_to_pes_19_out_bits = PE_349_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_37_io_to_pes_20_out_valid = PE_350_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_37_io_to_pes_20_out_bits = PE_350_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_37_io_to_mem_valid = MemController_37_io_rd_data_valid; // @[pe.scala 312:29]
  assign PENetwork_37_io_to_mem_bits = MemController_37_io_rd_data_bits; // @[pe.scala 312:29]
  assign PENetwork_38_io_to_pes_0_out_valid = PE_352_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_38_io_to_pes_0_out_bits = PE_352_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_38_io_to_pes_1_out_valid = PE_353_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_38_io_to_pes_1_out_bits = PE_353_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_38_io_to_pes_2_out_valid = PE_354_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_38_io_to_pes_2_out_bits = PE_354_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_38_io_to_pes_3_out_valid = PE_355_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_38_io_to_pes_3_out_bits = PE_355_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_38_io_to_pes_4_out_valid = PE_356_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_38_io_to_pes_4_out_bits = PE_356_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_38_io_to_pes_5_out_valid = PE_357_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_38_io_to_pes_5_out_bits = PE_357_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_38_io_to_pes_6_out_valid = PE_358_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_38_io_to_pes_6_out_bits = PE_358_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_38_io_to_pes_7_out_valid = PE_359_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_38_io_to_pes_7_out_bits = PE_359_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_38_io_to_pes_8_out_valid = PE_360_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_38_io_to_pes_8_out_bits = PE_360_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_38_io_to_pes_9_out_valid = PE_361_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_38_io_to_pes_9_out_bits = PE_361_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_38_io_to_pes_10_out_valid = PE_362_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_38_io_to_pes_10_out_bits = PE_362_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_38_io_to_pes_11_out_valid = PE_363_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_38_io_to_pes_11_out_bits = PE_363_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_38_io_to_pes_12_out_valid = PE_364_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_38_io_to_pes_12_out_bits = PE_364_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_38_io_to_pes_13_out_valid = PE_365_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_38_io_to_pes_13_out_bits = PE_365_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_38_io_to_pes_14_out_valid = PE_366_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_38_io_to_pes_14_out_bits = PE_366_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_38_io_to_pes_15_out_valid = PE_367_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_38_io_to_pes_15_out_bits = PE_367_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_38_io_to_pes_16_out_valid = PE_368_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_38_io_to_pes_16_out_bits = PE_368_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_38_io_to_pes_17_out_valid = PE_369_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_38_io_to_pes_17_out_bits = PE_369_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_38_io_to_pes_18_out_valid = PE_370_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_38_io_to_pes_18_out_bits = PE_370_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_38_io_to_pes_19_out_valid = PE_371_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_38_io_to_pes_19_out_bits = PE_371_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_38_io_to_pes_20_out_valid = PE_372_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_38_io_to_pes_20_out_bits = PE_372_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_38_io_to_mem_valid = MemController_38_io_rd_data_valid; // @[pe.scala 312:29]
  assign PENetwork_38_io_to_mem_bits = MemController_38_io_rd_data_bits; // @[pe.scala 312:29]
  assign PENetwork_39_io_to_pes_0_out_valid = PE_374_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_39_io_to_pes_0_out_bits = PE_374_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_39_io_to_pes_1_out_valid = PE_375_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_39_io_to_pes_1_out_bits = PE_375_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_39_io_to_pes_2_out_valid = PE_376_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_39_io_to_pes_2_out_bits = PE_376_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_39_io_to_pes_3_out_valid = PE_377_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_39_io_to_pes_3_out_bits = PE_377_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_39_io_to_pes_4_out_valid = PE_378_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_39_io_to_pes_4_out_bits = PE_378_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_39_io_to_pes_5_out_valid = PE_379_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_39_io_to_pes_5_out_bits = PE_379_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_39_io_to_pes_6_out_valid = PE_380_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_39_io_to_pes_6_out_bits = PE_380_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_39_io_to_pes_7_out_valid = PE_381_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_39_io_to_pes_7_out_bits = PE_381_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_39_io_to_pes_8_out_valid = PE_382_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_39_io_to_pes_8_out_bits = PE_382_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_39_io_to_pes_9_out_valid = PE_383_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_39_io_to_pes_9_out_bits = PE_383_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_39_io_to_pes_10_out_valid = PE_384_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_39_io_to_pes_10_out_bits = PE_384_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_39_io_to_pes_11_out_valid = PE_385_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_39_io_to_pes_11_out_bits = PE_385_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_39_io_to_pes_12_out_valid = PE_386_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_39_io_to_pes_12_out_bits = PE_386_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_39_io_to_pes_13_out_valid = PE_387_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_39_io_to_pes_13_out_bits = PE_387_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_39_io_to_pes_14_out_valid = PE_388_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_39_io_to_pes_14_out_bits = PE_388_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_39_io_to_pes_15_out_valid = PE_389_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_39_io_to_pes_15_out_bits = PE_389_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_39_io_to_pes_16_out_valid = PE_390_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_39_io_to_pes_16_out_bits = PE_390_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_39_io_to_pes_17_out_valid = PE_391_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_39_io_to_pes_17_out_bits = PE_391_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_39_io_to_pes_18_out_valid = PE_392_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_39_io_to_pes_18_out_bits = PE_392_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_39_io_to_pes_19_out_valid = PE_393_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_39_io_to_pes_19_out_bits = PE_393_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_39_io_to_pes_20_out_valid = PE_394_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_39_io_to_pes_20_out_bits = PE_394_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_39_io_to_mem_valid = MemController_39_io_rd_data_valid; // @[pe.scala 312:29]
  assign PENetwork_39_io_to_mem_bits = MemController_39_io_rd_data_bits; // @[pe.scala 312:29]
  assign PENetwork_40_io_to_pes_0_out_valid = PE_396_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_40_io_to_pes_0_out_bits = PE_396_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_40_io_to_pes_1_out_valid = PE_397_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_40_io_to_pes_1_out_bits = PE_397_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_40_io_to_pes_2_out_valid = PE_398_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_40_io_to_pes_2_out_bits = PE_398_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_40_io_to_pes_3_out_valid = PE_399_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_40_io_to_pes_3_out_bits = PE_399_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_40_io_to_pes_4_out_valid = PE_400_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_40_io_to_pes_4_out_bits = PE_400_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_40_io_to_pes_5_out_valid = PE_401_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_40_io_to_pes_5_out_bits = PE_401_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_40_io_to_pes_6_out_valid = PE_402_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_40_io_to_pes_6_out_bits = PE_402_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_40_io_to_pes_7_out_valid = PE_403_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_40_io_to_pes_7_out_bits = PE_403_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_40_io_to_pes_8_out_valid = PE_404_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_40_io_to_pes_8_out_bits = PE_404_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_40_io_to_pes_9_out_valid = PE_405_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_40_io_to_pes_9_out_bits = PE_405_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_40_io_to_pes_10_out_valid = PE_406_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_40_io_to_pes_10_out_bits = PE_406_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_40_io_to_pes_11_out_valid = PE_407_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_40_io_to_pes_11_out_bits = PE_407_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_40_io_to_pes_12_out_valid = PE_408_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_40_io_to_pes_12_out_bits = PE_408_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_40_io_to_pes_13_out_valid = PE_409_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_40_io_to_pes_13_out_bits = PE_409_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_40_io_to_pes_14_out_valid = PE_410_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_40_io_to_pes_14_out_bits = PE_410_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_40_io_to_pes_15_out_valid = PE_411_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_40_io_to_pes_15_out_bits = PE_411_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_40_io_to_pes_16_out_valid = PE_412_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_40_io_to_pes_16_out_bits = PE_412_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_40_io_to_pes_17_out_valid = PE_413_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_40_io_to_pes_17_out_bits = PE_413_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_40_io_to_pes_18_out_valid = PE_414_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_40_io_to_pes_18_out_bits = PE_414_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_40_io_to_pes_19_out_valid = PE_415_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_40_io_to_pes_19_out_bits = PE_415_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_40_io_to_pes_20_out_valid = PE_416_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_40_io_to_pes_20_out_bits = PE_416_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_40_io_to_mem_valid = MemController_40_io_rd_data_valid; // @[pe.scala 312:29]
  assign PENetwork_40_io_to_mem_bits = MemController_40_io_rd_data_bits; // @[pe.scala 312:29]
  assign PENetwork_41_io_to_pes_0_out_valid = PE_418_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_41_io_to_pes_0_out_bits = PE_418_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_41_io_to_pes_1_out_valid = PE_419_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_41_io_to_pes_1_out_bits = PE_419_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_41_io_to_pes_2_out_valid = PE_420_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_41_io_to_pes_2_out_bits = PE_420_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_41_io_to_pes_3_out_valid = PE_421_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_41_io_to_pes_3_out_bits = PE_421_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_41_io_to_pes_4_out_valid = PE_422_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_41_io_to_pes_4_out_bits = PE_422_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_41_io_to_pes_5_out_valid = PE_423_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_41_io_to_pes_5_out_bits = PE_423_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_41_io_to_pes_6_out_valid = PE_424_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_41_io_to_pes_6_out_bits = PE_424_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_41_io_to_pes_7_out_valid = PE_425_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_41_io_to_pes_7_out_bits = PE_425_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_41_io_to_pes_8_out_valid = PE_426_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_41_io_to_pes_8_out_bits = PE_426_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_41_io_to_pes_9_out_valid = PE_427_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_41_io_to_pes_9_out_bits = PE_427_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_41_io_to_pes_10_out_valid = PE_428_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_41_io_to_pes_10_out_bits = PE_428_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_41_io_to_pes_11_out_valid = PE_429_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_41_io_to_pes_11_out_bits = PE_429_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_41_io_to_pes_12_out_valid = PE_430_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_41_io_to_pes_12_out_bits = PE_430_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_41_io_to_pes_13_out_valid = PE_431_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_41_io_to_pes_13_out_bits = PE_431_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_41_io_to_pes_14_out_valid = PE_432_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_41_io_to_pes_14_out_bits = PE_432_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_41_io_to_pes_15_out_valid = PE_433_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_41_io_to_pes_15_out_bits = PE_433_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_41_io_to_pes_16_out_valid = PE_434_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_41_io_to_pes_16_out_bits = PE_434_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_41_io_to_pes_17_out_valid = PE_435_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_41_io_to_pes_17_out_bits = PE_435_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_41_io_to_pes_18_out_valid = PE_436_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_41_io_to_pes_18_out_bits = PE_436_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_41_io_to_pes_19_out_valid = PE_437_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_41_io_to_pes_19_out_bits = PE_437_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_41_io_to_pes_20_out_valid = PE_438_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_41_io_to_pes_20_out_bits = PE_438_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_41_io_to_mem_valid = MemController_41_io_rd_data_valid; // @[pe.scala 312:29]
  assign PENetwork_41_io_to_mem_bits = MemController_41_io_rd_data_bits; // @[pe.scala 312:29]
  assign PENetwork_42_io_to_pes_0_out_valid = PE_440_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_42_io_to_pes_0_out_bits = PE_440_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_42_io_to_pes_1_out_valid = PE_441_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_42_io_to_pes_1_out_bits = PE_441_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_42_io_to_pes_2_out_valid = PE_442_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_42_io_to_pes_2_out_bits = PE_442_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_42_io_to_pes_3_out_valid = PE_443_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_42_io_to_pes_3_out_bits = PE_443_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_42_io_to_pes_4_out_valid = PE_444_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_42_io_to_pes_4_out_bits = PE_444_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_42_io_to_pes_5_out_valid = PE_445_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_42_io_to_pes_5_out_bits = PE_445_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_42_io_to_pes_6_out_valid = PE_446_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_42_io_to_pes_6_out_bits = PE_446_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_42_io_to_pes_7_out_valid = PE_447_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_42_io_to_pes_7_out_bits = PE_447_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_42_io_to_pes_8_out_valid = PE_448_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_42_io_to_pes_8_out_bits = PE_448_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_42_io_to_pes_9_out_valid = PE_449_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_42_io_to_pes_9_out_bits = PE_449_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_42_io_to_pes_10_out_valid = PE_450_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_42_io_to_pes_10_out_bits = PE_450_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_42_io_to_pes_11_out_valid = PE_451_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_42_io_to_pes_11_out_bits = PE_451_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_42_io_to_pes_12_out_valid = PE_452_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_42_io_to_pes_12_out_bits = PE_452_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_42_io_to_pes_13_out_valid = PE_453_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_42_io_to_pes_13_out_bits = PE_453_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_42_io_to_pes_14_out_valid = PE_454_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_42_io_to_pes_14_out_bits = PE_454_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_42_io_to_pes_15_out_valid = PE_455_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_42_io_to_pes_15_out_bits = PE_455_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_42_io_to_pes_16_out_valid = PE_456_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_42_io_to_pes_16_out_bits = PE_456_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_42_io_to_pes_17_out_valid = PE_457_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_42_io_to_pes_17_out_bits = PE_457_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_42_io_to_pes_18_out_valid = PE_458_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_42_io_to_pes_18_out_bits = PE_458_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_42_io_to_pes_19_out_valid = PE_459_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_42_io_to_pes_19_out_bits = PE_459_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_42_io_to_pes_20_out_valid = PE_460_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_42_io_to_pes_20_out_bits = PE_460_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_42_io_to_mem_valid = MemController_42_io_rd_data_valid; // @[pe.scala 312:29]
  assign PENetwork_42_io_to_mem_bits = MemController_42_io_rd_data_bits; // @[pe.scala 312:29]
  assign PENetwork_43_io_to_pes_0_out_valid = PE_462_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_43_io_to_pes_0_out_bits = PE_462_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_43_io_to_pes_1_out_valid = PE_463_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_43_io_to_pes_1_out_bits = PE_463_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_43_io_to_pes_2_out_valid = PE_464_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_43_io_to_pes_2_out_bits = PE_464_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_43_io_to_pes_3_out_valid = PE_465_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_43_io_to_pes_3_out_bits = PE_465_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_43_io_to_pes_4_out_valid = PE_466_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_43_io_to_pes_4_out_bits = PE_466_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_43_io_to_pes_5_out_valid = PE_467_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_43_io_to_pes_5_out_bits = PE_467_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_43_io_to_pes_6_out_valid = PE_468_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_43_io_to_pes_6_out_bits = PE_468_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_43_io_to_pes_7_out_valid = PE_469_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_43_io_to_pes_7_out_bits = PE_469_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_43_io_to_pes_8_out_valid = PE_470_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_43_io_to_pes_8_out_bits = PE_470_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_43_io_to_pes_9_out_valid = PE_471_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_43_io_to_pes_9_out_bits = PE_471_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_43_io_to_pes_10_out_valid = PE_472_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_43_io_to_pes_10_out_bits = PE_472_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_43_io_to_pes_11_out_valid = PE_473_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_43_io_to_pes_11_out_bits = PE_473_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_43_io_to_pes_12_out_valid = PE_474_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_43_io_to_pes_12_out_bits = PE_474_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_43_io_to_pes_13_out_valid = PE_475_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_43_io_to_pes_13_out_bits = PE_475_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_43_io_to_pes_14_out_valid = PE_476_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_43_io_to_pes_14_out_bits = PE_476_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_43_io_to_pes_15_out_valid = PE_477_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_43_io_to_pes_15_out_bits = PE_477_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_43_io_to_pes_16_out_valid = PE_478_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_43_io_to_pes_16_out_bits = PE_478_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_43_io_to_pes_17_out_valid = PE_479_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_43_io_to_pes_17_out_bits = PE_479_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_43_io_to_pes_18_out_valid = PE_480_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_43_io_to_pes_18_out_bits = PE_480_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_43_io_to_pes_19_out_valid = PE_481_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_43_io_to_pes_19_out_bits = PE_481_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_43_io_to_pes_20_out_valid = PE_482_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_43_io_to_pes_20_out_bits = PE_482_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_43_io_to_mem_valid = MemController_43_io_rd_data_valid; // @[pe.scala 312:29]
  assign PENetwork_43_io_to_mem_bits = MemController_43_io_rd_data_bits; // @[pe.scala 312:29]
  assign PENetwork_44_io_to_pes_0_out_valid = PE_484_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_44_io_to_pes_0_out_bits = PE_484_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_44_io_to_pes_1_out_valid = PE_485_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_44_io_to_pes_1_out_bits = PE_485_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_44_io_to_pes_2_out_valid = PE_486_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_44_io_to_pes_2_out_bits = PE_486_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_44_io_to_pes_3_out_valid = PE_487_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_44_io_to_pes_3_out_bits = PE_487_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_44_io_to_pes_4_out_valid = PE_488_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_44_io_to_pes_4_out_bits = PE_488_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_44_io_to_pes_5_out_valid = PE_489_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_44_io_to_pes_5_out_bits = PE_489_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_44_io_to_pes_6_out_valid = PE_490_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_44_io_to_pes_6_out_bits = PE_490_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_44_io_to_pes_7_out_valid = PE_491_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_44_io_to_pes_7_out_bits = PE_491_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_44_io_to_pes_8_out_valid = PE_492_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_44_io_to_pes_8_out_bits = PE_492_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_44_io_to_pes_9_out_valid = PE_493_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_44_io_to_pes_9_out_bits = PE_493_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_44_io_to_pes_10_out_valid = PE_494_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_44_io_to_pes_10_out_bits = PE_494_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_44_io_to_pes_11_out_valid = PE_495_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_44_io_to_pes_11_out_bits = PE_495_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_44_io_to_pes_12_out_valid = PE_496_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_44_io_to_pes_12_out_bits = PE_496_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_44_io_to_pes_13_out_valid = PE_497_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_44_io_to_pes_13_out_bits = PE_497_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_44_io_to_pes_14_out_valid = PE_498_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_44_io_to_pes_14_out_bits = PE_498_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_44_io_to_pes_15_out_valid = PE_499_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_44_io_to_pes_15_out_bits = PE_499_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_44_io_to_pes_16_out_valid = PE_500_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_44_io_to_pes_16_out_bits = PE_500_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_44_io_to_pes_17_out_valid = PE_501_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_44_io_to_pes_17_out_bits = PE_501_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_44_io_to_pes_18_out_valid = PE_502_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_44_io_to_pes_18_out_bits = PE_502_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_44_io_to_pes_19_out_valid = PE_503_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_44_io_to_pes_19_out_bits = PE_503_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_44_io_to_pes_20_out_valid = PE_504_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_44_io_to_pes_20_out_bits = PE_504_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_44_io_to_mem_valid = MemController_44_io_rd_data_valid; // @[pe.scala 312:29]
  assign PENetwork_44_io_to_mem_bits = MemController_44_io_rd_data_bits; // @[pe.scala 312:29]
  assign PENetwork_45_io_to_pes_0_out_valid = PE_506_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_45_io_to_pes_0_out_bits = PE_506_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_45_io_to_pes_1_out_valid = PE_507_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_45_io_to_pes_1_out_bits = PE_507_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_45_io_to_pes_2_out_valid = PE_508_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_45_io_to_pes_2_out_bits = PE_508_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_45_io_to_pes_3_out_valid = PE_509_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_45_io_to_pes_3_out_bits = PE_509_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_45_io_to_pes_4_out_valid = PE_510_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_45_io_to_pes_4_out_bits = PE_510_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_45_io_to_pes_5_out_valid = PE_511_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_45_io_to_pes_5_out_bits = PE_511_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_45_io_to_pes_6_out_valid = PE_512_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_45_io_to_pes_6_out_bits = PE_512_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_45_io_to_pes_7_out_valid = PE_513_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_45_io_to_pes_7_out_bits = PE_513_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_45_io_to_pes_8_out_valid = PE_514_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_45_io_to_pes_8_out_bits = PE_514_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_45_io_to_pes_9_out_valid = PE_515_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_45_io_to_pes_9_out_bits = PE_515_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_45_io_to_pes_10_out_valid = PE_516_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_45_io_to_pes_10_out_bits = PE_516_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_45_io_to_pes_11_out_valid = PE_517_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_45_io_to_pes_11_out_bits = PE_517_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_45_io_to_pes_12_out_valid = PE_518_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_45_io_to_pes_12_out_bits = PE_518_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_45_io_to_pes_13_out_valid = PE_519_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_45_io_to_pes_13_out_bits = PE_519_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_45_io_to_pes_14_out_valid = PE_520_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_45_io_to_pes_14_out_bits = PE_520_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_45_io_to_pes_15_out_valid = PE_521_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_45_io_to_pes_15_out_bits = PE_521_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_45_io_to_pes_16_out_valid = PE_522_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_45_io_to_pes_16_out_bits = PE_522_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_45_io_to_pes_17_out_valid = PE_523_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_45_io_to_pes_17_out_bits = PE_523_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_45_io_to_pes_18_out_valid = PE_524_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_45_io_to_pes_18_out_bits = PE_524_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_45_io_to_pes_19_out_valid = PE_525_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_45_io_to_pes_19_out_bits = PE_525_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_45_io_to_pes_20_out_valid = PE_526_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_45_io_to_pes_20_out_bits = PE_526_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_45_io_to_mem_valid = MemController_45_io_rd_data_valid; // @[pe.scala 312:29]
  assign PENetwork_45_io_to_mem_bits = MemController_45_io_rd_data_bits; // @[pe.scala 312:29]
  assign PENetwork_46_io_to_pes_0_out_valid = PE_528_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_46_io_to_pes_0_out_bits = PE_528_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_46_io_to_pes_1_out_valid = PE_529_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_46_io_to_pes_1_out_bits = PE_529_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_46_io_to_pes_2_out_valid = PE_530_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_46_io_to_pes_2_out_bits = PE_530_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_46_io_to_pes_3_out_valid = PE_531_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_46_io_to_pes_3_out_bits = PE_531_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_46_io_to_pes_4_out_valid = PE_532_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_46_io_to_pes_4_out_bits = PE_532_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_46_io_to_pes_5_out_valid = PE_533_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_46_io_to_pes_5_out_bits = PE_533_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_46_io_to_pes_6_out_valid = PE_534_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_46_io_to_pes_6_out_bits = PE_534_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_46_io_to_pes_7_out_valid = PE_535_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_46_io_to_pes_7_out_bits = PE_535_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_46_io_to_pes_8_out_valid = PE_536_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_46_io_to_pes_8_out_bits = PE_536_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_46_io_to_pes_9_out_valid = PE_537_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_46_io_to_pes_9_out_bits = PE_537_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_46_io_to_pes_10_out_valid = PE_538_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_46_io_to_pes_10_out_bits = PE_538_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_46_io_to_pes_11_out_valid = PE_539_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_46_io_to_pes_11_out_bits = PE_539_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_46_io_to_pes_12_out_valid = PE_540_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_46_io_to_pes_12_out_bits = PE_540_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_46_io_to_pes_13_out_valid = PE_541_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_46_io_to_pes_13_out_bits = PE_541_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_46_io_to_pes_14_out_valid = PE_542_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_46_io_to_pes_14_out_bits = PE_542_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_46_io_to_pes_15_out_valid = PE_543_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_46_io_to_pes_15_out_bits = PE_543_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_46_io_to_pes_16_out_valid = PE_544_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_46_io_to_pes_16_out_bits = PE_544_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_46_io_to_pes_17_out_valid = PE_545_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_46_io_to_pes_17_out_bits = PE_545_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_46_io_to_pes_18_out_valid = PE_546_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_46_io_to_pes_18_out_bits = PE_546_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_46_io_to_pes_19_out_valid = PE_547_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_46_io_to_pes_19_out_bits = PE_547_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_46_io_to_pes_20_out_valid = PE_548_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_46_io_to_pes_20_out_bits = PE_548_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_46_io_to_mem_valid = MemController_46_io_rd_data_valid; // @[pe.scala 312:29]
  assign PENetwork_46_io_to_mem_bits = MemController_46_io_rd_data_bits; // @[pe.scala 312:29]
  assign PENetwork_47_io_to_pes_0_out_valid = PE_550_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_47_io_to_pes_0_out_bits = PE_550_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_47_io_to_pes_1_out_valid = PE_551_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_47_io_to_pes_1_out_bits = PE_551_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_47_io_to_pes_2_out_valid = PE_552_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_47_io_to_pes_2_out_bits = PE_552_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_47_io_to_pes_3_out_valid = PE_553_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_47_io_to_pes_3_out_bits = PE_553_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_47_io_to_pes_4_out_valid = PE_554_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_47_io_to_pes_4_out_bits = PE_554_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_47_io_to_pes_5_out_valid = PE_555_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_47_io_to_pes_5_out_bits = PE_555_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_47_io_to_pes_6_out_valid = PE_556_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_47_io_to_pes_6_out_bits = PE_556_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_47_io_to_pes_7_out_valid = PE_557_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_47_io_to_pes_7_out_bits = PE_557_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_47_io_to_pes_8_out_valid = PE_558_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_47_io_to_pes_8_out_bits = PE_558_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_47_io_to_pes_9_out_valid = PE_559_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_47_io_to_pes_9_out_bits = PE_559_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_47_io_to_pes_10_out_valid = PE_560_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_47_io_to_pes_10_out_bits = PE_560_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_47_io_to_pes_11_out_valid = PE_561_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_47_io_to_pes_11_out_bits = PE_561_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_47_io_to_pes_12_out_valid = PE_562_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_47_io_to_pes_12_out_bits = PE_562_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_47_io_to_pes_13_out_valid = PE_563_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_47_io_to_pes_13_out_bits = PE_563_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_47_io_to_pes_14_out_valid = PE_564_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_47_io_to_pes_14_out_bits = PE_564_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_47_io_to_pes_15_out_valid = PE_565_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_47_io_to_pes_15_out_bits = PE_565_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_47_io_to_pes_16_out_valid = PE_566_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_47_io_to_pes_16_out_bits = PE_566_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_47_io_to_pes_17_out_valid = PE_567_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_47_io_to_pes_17_out_bits = PE_567_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_47_io_to_pes_18_out_valid = PE_568_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_47_io_to_pes_18_out_bits = PE_568_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_47_io_to_pes_19_out_valid = PE_569_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_47_io_to_pes_19_out_bits = PE_569_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_47_io_to_pes_20_out_valid = PE_570_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_47_io_to_pes_20_out_bits = PE_570_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_47_io_to_mem_valid = MemController_47_io_rd_data_valid; // @[pe.scala 312:29]
  assign PENetwork_47_io_to_mem_bits = MemController_47_io_rd_data_bits; // @[pe.scala 312:29]
  assign PENetwork_48_io_to_pes_0_out_valid = PE_572_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_48_io_to_pes_0_out_bits = PE_572_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_48_io_to_pes_1_out_valid = PE_573_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_48_io_to_pes_1_out_bits = PE_573_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_48_io_to_pes_2_out_valid = PE_574_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_48_io_to_pes_2_out_bits = PE_574_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_48_io_to_pes_3_out_valid = PE_575_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_48_io_to_pes_3_out_bits = PE_575_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_48_io_to_pes_4_out_valid = PE_576_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_48_io_to_pes_4_out_bits = PE_576_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_48_io_to_pes_5_out_valid = PE_577_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_48_io_to_pes_5_out_bits = PE_577_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_48_io_to_pes_6_out_valid = PE_578_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_48_io_to_pes_6_out_bits = PE_578_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_48_io_to_pes_7_out_valid = PE_579_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_48_io_to_pes_7_out_bits = PE_579_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_48_io_to_pes_8_out_valid = PE_580_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_48_io_to_pes_8_out_bits = PE_580_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_48_io_to_pes_9_out_valid = PE_581_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_48_io_to_pes_9_out_bits = PE_581_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_48_io_to_pes_10_out_valid = PE_582_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_48_io_to_pes_10_out_bits = PE_582_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_48_io_to_pes_11_out_valid = PE_583_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_48_io_to_pes_11_out_bits = PE_583_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_48_io_to_pes_12_out_valid = PE_584_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_48_io_to_pes_12_out_bits = PE_584_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_48_io_to_pes_13_out_valid = PE_585_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_48_io_to_pes_13_out_bits = PE_585_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_48_io_to_pes_14_out_valid = PE_586_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_48_io_to_pes_14_out_bits = PE_586_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_48_io_to_pes_15_out_valid = PE_587_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_48_io_to_pes_15_out_bits = PE_587_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_48_io_to_pes_16_out_valid = PE_588_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_48_io_to_pes_16_out_bits = PE_588_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_48_io_to_pes_17_out_valid = PE_589_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_48_io_to_pes_17_out_bits = PE_589_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_48_io_to_pes_18_out_valid = PE_590_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_48_io_to_pes_18_out_bits = PE_590_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_48_io_to_pes_19_out_valid = PE_591_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_48_io_to_pes_19_out_bits = PE_591_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_48_io_to_pes_20_out_valid = PE_592_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_48_io_to_pes_20_out_bits = PE_592_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_48_io_to_mem_valid = MemController_48_io_rd_data_valid; // @[pe.scala 312:29]
  assign PENetwork_48_io_to_mem_bits = MemController_48_io_rd_data_bits; // @[pe.scala 312:29]
  assign PENetwork_49_io_to_pes_0_out_valid = PE_594_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_49_io_to_pes_0_out_bits = PE_594_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_49_io_to_pes_1_out_valid = PE_595_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_49_io_to_pes_1_out_bits = PE_595_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_49_io_to_pes_2_out_valid = PE_596_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_49_io_to_pes_2_out_bits = PE_596_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_49_io_to_pes_3_out_valid = PE_597_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_49_io_to_pes_3_out_bits = PE_597_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_49_io_to_pes_4_out_valid = PE_598_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_49_io_to_pes_4_out_bits = PE_598_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_49_io_to_pes_5_out_valid = PE_599_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_49_io_to_pes_5_out_bits = PE_599_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_49_io_to_pes_6_out_valid = PE_600_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_49_io_to_pes_6_out_bits = PE_600_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_49_io_to_pes_7_out_valid = PE_601_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_49_io_to_pes_7_out_bits = PE_601_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_49_io_to_pes_8_out_valid = PE_602_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_49_io_to_pes_8_out_bits = PE_602_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_49_io_to_pes_9_out_valid = PE_603_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_49_io_to_pes_9_out_bits = PE_603_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_49_io_to_pes_10_out_valid = PE_604_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_49_io_to_pes_10_out_bits = PE_604_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_49_io_to_pes_11_out_valid = PE_605_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_49_io_to_pes_11_out_bits = PE_605_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_49_io_to_pes_12_out_valid = PE_606_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_49_io_to_pes_12_out_bits = PE_606_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_49_io_to_pes_13_out_valid = PE_607_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_49_io_to_pes_13_out_bits = PE_607_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_49_io_to_pes_14_out_valid = PE_608_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_49_io_to_pes_14_out_bits = PE_608_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_49_io_to_pes_15_out_valid = PE_609_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_49_io_to_pes_15_out_bits = PE_609_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_49_io_to_pes_16_out_valid = PE_610_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_49_io_to_pes_16_out_bits = PE_610_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_49_io_to_pes_17_out_valid = PE_611_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_49_io_to_pes_17_out_bits = PE_611_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_49_io_to_pes_18_out_valid = PE_612_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_49_io_to_pes_18_out_bits = PE_612_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_49_io_to_pes_19_out_valid = PE_613_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_49_io_to_pes_19_out_bits = PE_613_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_49_io_to_pes_20_out_valid = PE_614_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_49_io_to_pes_20_out_bits = PE_614_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_49_io_to_mem_valid = MemController_49_io_rd_data_valid; // @[pe.scala 312:29]
  assign PENetwork_49_io_to_mem_bits = MemController_49_io_rd_data_bits; // @[pe.scala 312:29]
  assign PENetwork_50_io_to_pes_0_out_valid = PE_616_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_50_io_to_pes_0_out_bits = PE_616_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_50_io_to_pes_1_out_valid = PE_617_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_50_io_to_pes_1_out_bits = PE_617_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_50_io_to_pes_2_out_valid = PE_618_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_50_io_to_pes_2_out_bits = PE_618_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_50_io_to_pes_3_out_valid = PE_619_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_50_io_to_pes_3_out_bits = PE_619_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_50_io_to_pes_4_out_valid = PE_620_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_50_io_to_pes_4_out_bits = PE_620_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_50_io_to_pes_5_out_valid = PE_621_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_50_io_to_pes_5_out_bits = PE_621_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_50_io_to_pes_6_out_valid = PE_622_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_50_io_to_pes_6_out_bits = PE_622_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_50_io_to_pes_7_out_valid = PE_623_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_50_io_to_pes_7_out_bits = PE_623_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_50_io_to_pes_8_out_valid = PE_624_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_50_io_to_pes_8_out_bits = PE_624_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_50_io_to_pes_9_out_valid = PE_625_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_50_io_to_pes_9_out_bits = PE_625_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_50_io_to_pes_10_out_valid = PE_626_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_50_io_to_pes_10_out_bits = PE_626_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_50_io_to_pes_11_out_valid = PE_627_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_50_io_to_pes_11_out_bits = PE_627_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_50_io_to_pes_12_out_valid = PE_628_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_50_io_to_pes_12_out_bits = PE_628_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_50_io_to_pes_13_out_valid = PE_629_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_50_io_to_pes_13_out_bits = PE_629_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_50_io_to_pes_14_out_valid = PE_630_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_50_io_to_pes_14_out_bits = PE_630_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_50_io_to_pes_15_out_valid = PE_631_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_50_io_to_pes_15_out_bits = PE_631_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_50_io_to_pes_16_out_valid = PE_632_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_50_io_to_pes_16_out_bits = PE_632_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_50_io_to_pes_17_out_valid = PE_633_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_50_io_to_pes_17_out_bits = PE_633_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_50_io_to_pes_18_out_valid = PE_634_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_50_io_to_pes_18_out_bits = PE_634_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_50_io_to_pes_19_out_valid = PE_635_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_50_io_to_pes_19_out_bits = PE_635_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_50_io_to_pes_20_out_valid = PE_636_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_50_io_to_pes_20_out_bits = PE_636_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_50_io_to_mem_valid = MemController_50_io_rd_data_valid; // @[pe.scala 312:29]
  assign PENetwork_50_io_to_mem_bits = MemController_50_io_rd_data_bits; // @[pe.scala 312:29]
  assign PENetwork_51_io_to_pes_0_out_valid = PE_638_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_51_io_to_pes_0_out_bits = PE_638_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_51_io_to_pes_1_out_valid = PE_639_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_51_io_to_pes_1_out_bits = PE_639_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_51_io_to_pes_2_out_valid = PE_640_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_51_io_to_pes_2_out_bits = PE_640_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_51_io_to_pes_3_out_valid = PE_641_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_51_io_to_pes_3_out_bits = PE_641_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_51_io_to_pes_4_out_valid = PE_642_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_51_io_to_pes_4_out_bits = PE_642_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_51_io_to_pes_5_out_valid = PE_643_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_51_io_to_pes_5_out_bits = PE_643_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_51_io_to_pes_6_out_valid = PE_644_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_51_io_to_pes_6_out_bits = PE_644_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_51_io_to_pes_7_out_valid = PE_645_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_51_io_to_pes_7_out_bits = PE_645_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_51_io_to_pes_8_out_valid = PE_646_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_51_io_to_pes_8_out_bits = PE_646_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_51_io_to_pes_9_out_valid = PE_647_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_51_io_to_pes_9_out_bits = PE_647_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_51_io_to_pes_10_out_valid = PE_648_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_51_io_to_pes_10_out_bits = PE_648_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_51_io_to_pes_11_out_valid = PE_649_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_51_io_to_pes_11_out_bits = PE_649_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_51_io_to_pes_12_out_valid = PE_650_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_51_io_to_pes_12_out_bits = PE_650_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_51_io_to_pes_13_out_valid = PE_651_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_51_io_to_pes_13_out_bits = PE_651_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_51_io_to_pes_14_out_valid = PE_652_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_51_io_to_pes_14_out_bits = PE_652_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_51_io_to_pes_15_out_valid = PE_653_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_51_io_to_pes_15_out_bits = PE_653_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_51_io_to_pes_16_out_valid = PE_654_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_51_io_to_pes_16_out_bits = PE_654_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_51_io_to_pes_17_out_valid = PE_655_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_51_io_to_pes_17_out_bits = PE_655_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_51_io_to_pes_18_out_valid = PE_656_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_51_io_to_pes_18_out_bits = PE_656_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_51_io_to_pes_19_out_valid = PE_657_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_51_io_to_pes_19_out_bits = PE_657_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_51_io_to_pes_20_out_valid = PE_658_io_data_1_out_valid; // @[pe.scala 263:36]
  assign PENetwork_51_io_to_pes_20_out_bits = PE_658_io_data_1_out_bits; // @[pe.scala 263:36]
  assign PENetwork_51_io_to_mem_valid = MemController_51_io_rd_data_valid; // @[pe.scala 312:29]
  assign PENetwork_51_io_to_mem_bits = MemController_51_io_rd_data_bits; // @[pe.scala 312:29]
  assign PENetwork_52_clock = clock;
  assign PENetwork_52_reset = reset;
  assign PENetwork_52_io_to_pes_0_out_valid = PE_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_52_io_to_pes_0_out_bits = PE_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_52_io_to_pes_1_out_valid = PE_1_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_52_io_to_pes_1_out_bits = PE_1_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_52_io_to_pes_2_out_valid = PE_2_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_52_io_to_pes_2_out_bits = PE_2_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_52_io_to_pes_3_out_valid = PE_3_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_52_io_to_pes_3_out_bits = PE_3_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_52_io_to_pes_4_out_valid = PE_4_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_52_io_to_pes_4_out_bits = PE_4_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_52_io_to_pes_5_out_valid = PE_5_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_52_io_to_pes_5_out_bits = PE_5_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_52_io_to_pes_6_out_valid = PE_6_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_52_io_to_pes_6_out_bits = PE_6_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_52_io_to_pes_7_out_valid = PE_7_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_52_io_to_pes_7_out_bits = PE_7_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_52_io_to_pes_8_out_valid = PE_8_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_52_io_to_pes_8_out_bits = PE_8_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_52_io_to_pes_9_out_valid = PE_9_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_52_io_to_pes_9_out_bits = PE_9_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_52_io_to_pes_10_out_valid = PE_10_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_52_io_to_pes_10_out_bits = PE_10_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_52_io_to_pes_11_out_valid = PE_11_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_52_io_to_pes_11_out_bits = PE_11_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_52_io_to_pes_12_out_valid = PE_12_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_52_io_to_pes_12_out_bits = PE_12_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_52_io_to_pes_13_out_valid = PE_13_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_52_io_to_pes_13_out_bits = PE_13_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_52_io_to_pes_14_out_valid = PE_14_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_52_io_to_pes_14_out_bits = PE_14_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_52_io_to_pes_15_out_valid = PE_15_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_52_io_to_pes_15_out_bits = PE_15_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_52_io_to_pes_16_out_valid = PE_16_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_52_io_to_pes_16_out_bits = PE_16_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_52_io_to_pes_17_out_valid = PE_17_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_52_io_to_pes_17_out_bits = PE_17_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_52_io_to_pes_18_out_valid = PE_18_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_52_io_to_pes_18_out_bits = PE_18_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_52_io_to_pes_19_out_valid = PE_19_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_52_io_to_pes_19_out_bits = PE_19_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_52_io_to_pes_20_out_valid = PE_20_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_52_io_to_pes_20_out_bits = PE_20_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_52_io_to_pes_21_out_valid = PE_21_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_52_io_to_pes_21_out_bits = PE_21_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_52_io_sig_stat2trans = MultiDimTime_io_index_1 == 16'h0; // @[pe.scala 278:43]
  assign PENetwork_53_clock = clock;
  assign PENetwork_53_reset = reset;
  assign PENetwork_53_io_to_pes_0_out_valid = PE_22_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_53_io_to_pes_0_out_bits = PE_22_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_53_io_to_pes_1_out_valid = PE_23_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_53_io_to_pes_1_out_bits = PE_23_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_53_io_to_pes_2_out_valid = PE_24_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_53_io_to_pes_2_out_bits = PE_24_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_53_io_to_pes_3_out_valid = PE_25_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_53_io_to_pes_3_out_bits = PE_25_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_53_io_to_pes_4_out_valid = PE_26_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_53_io_to_pes_4_out_bits = PE_26_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_53_io_to_pes_5_out_valid = PE_27_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_53_io_to_pes_5_out_bits = PE_27_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_53_io_to_pes_6_out_valid = PE_28_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_53_io_to_pes_6_out_bits = PE_28_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_53_io_to_pes_7_out_valid = PE_29_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_53_io_to_pes_7_out_bits = PE_29_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_53_io_to_pes_8_out_valid = PE_30_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_53_io_to_pes_8_out_bits = PE_30_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_53_io_to_pes_9_out_valid = PE_31_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_53_io_to_pes_9_out_bits = PE_31_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_53_io_to_pes_10_out_valid = PE_32_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_53_io_to_pes_10_out_bits = PE_32_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_53_io_to_pes_11_out_valid = PE_33_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_53_io_to_pes_11_out_bits = PE_33_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_53_io_to_pes_12_out_valid = PE_34_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_53_io_to_pes_12_out_bits = PE_34_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_53_io_to_pes_13_out_valid = PE_35_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_53_io_to_pes_13_out_bits = PE_35_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_53_io_to_pes_14_out_valid = PE_36_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_53_io_to_pes_14_out_bits = PE_36_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_53_io_to_pes_15_out_valid = PE_37_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_53_io_to_pes_15_out_bits = PE_37_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_53_io_to_pes_16_out_valid = PE_38_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_53_io_to_pes_16_out_bits = PE_38_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_53_io_to_pes_17_out_valid = PE_39_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_53_io_to_pes_17_out_bits = PE_39_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_53_io_to_pes_18_out_valid = PE_40_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_53_io_to_pes_18_out_bits = PE_40_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_53_io_to_pes_19_out_valid = PE_41_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_53_io_to_pes_19_out_bits = PE_41_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_53_io_to_pes_20_out_valid = PE_42_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_53_io_to_pes_20_out_bits = PE_42_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_53_io_to_pes_21_out_valid = PE_43_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_53_io_to_pes_21_out_bits = PE_43_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_53_io_sig_stat2trans = MultiDimTime_io_index_1 == 16'h0; // @[pe.scala 278:43]
  assign PENetwork_54_clock = clock;
  assign PENetwork_54_reset = reset;
  assign PENetwork_54_io_to_pes_0_out_valid = PE_44_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_54_io_to_pes_0_out_bits = PE_44_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_54_io_to_pes_1_out_valid = PE_45_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_54_io_to_pes_1_out_bits = PE_45_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_54_io_to_pes_2_out_valid = PE_46_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_54_io_to_pes_2_out_bits = PE_46_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_54_io_to_pes_3_out_valid = PE_47_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_54_io_to_pes_3_out_bits = PE_47_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_54_io_to_pes_4_out_valid = PE_48_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_54_io_to_pes_4_out_bits = PE_48_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_54_io_to_pes_5_out_valid = PE_49_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_54_io_to_pes_5_out_bits = PE_49_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_54_io_to_pes_6_out_valid = PE_50_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_54_io_to_pes_6_out_bits = PE_50_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_54_io_to_pes_7_out_valid = PE_51_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_54_io_to_pes_7_out_bits = PE_51_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_54_io_to_pes_8_out_valid = PE_52_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_54_io_to_pes_8_out_bits = PE_52_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_54_io_to_pes_9_out_valid = PE_53_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_54_io_to_pes_9_out_bits = PE_53_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_54_io_to_pes_10_out_valid = PE_54_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_54_io_to_pes_10_out_bits = PE_54_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_54_io_to_pes_11_out_valid = PE_55_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_54_io_to_pes_11_out_bits = PE_55_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_54_io_to_pes_12_out_valid = PE_56_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_54_io_to_pes_12_out_bits = PE_56_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_54_io_to_pes_13_out_valid = PE_57_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_54_io_to_pes_13_out_bits = PE_57_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_54_io_to_pes_14_out_valid = PE_58_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_54_io_to_pes_14_out_bits = PE_58_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_54_io_to_pes_15_out_valid = PE_59_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_54_io_to_pes_15_out_bits = PE_59_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_54_io_to_pes_16_out_valid = PE_60_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_54_io_to_pes_16_out_bits = PE_60_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_54_io_to_pes_17_out_valid = PE_61_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_54_io_to_pes_17_out_bits = PE_61_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_54_io_to_pes_18_out_valid = PE_62_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_54_io_to_pes_18_out_bits = PE_62_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_54_io_to_pes_19_out_valid = PE_63_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_54_io_to_pes_19_out_bits = PE_63_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_54_io_to_pes_20_out_valid = PE_64_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_54_io_to_pes_20_out_bits = PE_64_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_54_io_to_pes_21_out_valid = PE_65_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_54_io_to_pes_21_out_bits = PE_65_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_54_io_sig_stat2trans = MultiDimTime_io_index_1 == 16'h0; // @[pe.scala 278:43]
  assign PENetwork_55_clock = clock;
  assign PENetwork_55_reset = reset;
  assign PENetwork_55_io_to_pes_0_out_valid = PE_66_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_55_io_to_pes_0_out_bits = PE_66_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_55_io_to_pes_1_out_valid = PE_67_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_55_io_to_pes_1_out_bits = PE_67_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_55_io_to_pes_2_out_valid = PE_68_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_55_io_to_pes_2_out_bits = PE_68_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_55_io_to_pes_3_out_valid = PE_69_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_55_io_to_pes_3_out_bits = PE_69_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_55_io_to_pes_4_out_valid = PE_70_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_55_io_to_pes_4_out_bits = PE_70_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_55_io_to_pes_5_out_valid = PE_71_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_55_io_to_pes_5_out_bits = PE_71_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_55_io_to_pes_6_out_valid = PE_72_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_55_io_to_pes_6_out_bits = PE_72_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_55_io_to_pes_7_out_valid = PE_73_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_55_io_to_pes_7_out_bits = PE_73_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_55_io_to_pes_8_out_valid = PE_74_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_55_io_to_pes_8_out_bits = PE_74_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_55_io_to_pes_9_out_valid = PE_75_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_55_io_to_pes_9_out_bits = PE_75_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_55_io_to_pes_10_out_valid = PE_76_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_55_io_to_pes_10_out_bits = PE_76_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_55_io_to_pes_11_out_valid = PE_77_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_55_io_to_pes_11_out_bits = PE_77_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_55_io_to_pes_12_out_valid = PE_78_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_55_io_to_pes_12_out_bits = PE_78_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_55_io_to_pes_13_out_valid = PE_79_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_55_io_to_pes_13_out_bits = PE_79_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_55_io_to_pes_14_out_valid = PE_80_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_55_io_to_pes_14_out_bits = PE_80_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_55_io_to_pes_15_out_valid = PE_81_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_55_io_to_pes_15_out_bits = PE_81_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_55_io_to_pes_16_out_valid = PE_82_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_55_io_to_pes_16_out_bits = PE_82_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_55_io_to_pes_17_out_valid = PE_83_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_55_io_to_pes_17_out_bits = PE_83_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_55_io_to_pes_18_out_valid = PE_84_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_55_io_to_pes_18_out_bits = PE_84_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_55_io_to_pes_19_out_valid = PE_85_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_55_io_to_pes_19_out_bits = PE_85_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_55_io_to_pes_20_out_valid = PE_86_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_55_io_to_pes_20_out_bits = PE_86_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_55_io_to_pes_21_out_valid = PE_87_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_55_io_to_pes_21_out_bits = PE_87_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_55_io_sig_stat2trans = MultiDimTime_io_index_1 == 16'h0; // @[pe.scala 278:43]
  assign PENetwork_56_clock = clock;
  assign PENetwork_56_reset = reset;
  assign PENetwork_56_io_to_pes_0_out_valid = PE_88_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_56_io_to_pes_0_out_bits = PE_88_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_56_io_to_pes_1_out_valid = PE_89_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_56_io_to_pes_1_out_bits = PE_89_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_56_io_to_pes_2_out_valid = PE_90_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_56_io_to_pes_2_out_bits = PE_90_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_56_io_to_pes_3_out_valid = PE_91_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_56_io_to_pes_3_out_bits = PE_91_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_56_io_to_pes_4_out_valid = PE_92_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_56_io_to_pes_4_out_bits = PE_92_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_56_io_to_pes_5_out_valid = PE_93_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_56_io_to_pes_5_out_bits = PE_93_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_56_io_to_pes_6_out_valid = PE_94_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_56_io_to_pes_6_out_bits = PE_94_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_56_io_to_pes_7_out_valid = PE_95_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_56_io_to_pes_7_out_bits = PE_95_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_56_io_to_pes_8_out_valid = PE_96_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_56_io_to_pes_8_out_bits = PE_96_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_56_io_to_pes_9_out_valid = PE_97_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_56_io_to_pes_9_out_bits = PE_97_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_56_io_to_pes_10_out_valid = PE_98_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_56_io_to_pes_10_out_bits = PE_98_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_56_io_to_pes_11_out_valid = PE_99_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_56_io_to_pes_11_out_bits = PE_99_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_56_io_to_pes_12_out_valid = PE_100_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_56_io_to_pes_12_out_bits = PE_100_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_56_io_to_pes_13_out_valid = PE_101_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_56_io_to_pes_13_out_bits = PE_101_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_56_io_to_pes_14_out_valid = PE_102_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_56_io_to_pes_14_out_bits = PE_102_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_56_io_to_pes_15_out_valid = PE_103_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_56_io_to_pes_15_out_bits = PE_103_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_56_io_to_pes_16_out_valid = PE_104_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_56_io_to_pes_16_out_bits = PE_104_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_56_io_to_pes_17_out_valid = PE_105_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_56_io_to_pes_17_out_bits = PE_105_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_56_io_to_pes_18_out_valid = PE_106_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_56_io_to_pes_18_out_bits = PE_106_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_56_io_to_pes_19_out_valid = PE_107_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_56_io_to_pes_19_out_bits = PE_107_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_56_io_to_pes_20_out_valid = PE_108_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_56_io_to_pes_20_out_bits = PE_108_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_56_io_to_pes_21_out_valid = PE_109_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_56_io_to_pes_21_out_bits = PE_109_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_56_io_sig_stat2trans = MultiDimTime_io_index_1 == 16'h0; // @[pe.scala 278:43]
  assign PENetwork_57_clock = clock;
  assign PENetwork_57_reset = reset;
  assign PENetwork_57_io_to_pes_0_out_valid = PE_110_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_57_io_to_pes_0_out_bits = PE_110_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_57_io_to_pes_1_out_valid = PE_111_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_57_io_to_pes_1_out_bits = PE_111_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_57_io_to_pes_2_out_valid = PE_112_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_57_io_to_pes_2_out_bits = PE_112_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_57_io_to_pes_3_out_valid = PE_113_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_57_io_to_pes_3_out_bits = PE_113_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_57_io_to_pes_4_out_valid = PE_114_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_57_io_to_pes_4_out_bits = PE_114_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_57_io_to_pes_5_out_valid = PE_115_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_57_io_to_pes_5_out_bits = PE_115_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_57_io_to_pes_6_out_valid = PE_116_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_57_io_to_pes_6_out_bits = PE_116_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_57_io_to_pes_7_out_valid = PE_117_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_57_io_to_pes_7_out_bits = PE_117_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_57_io_to_pes_8_out_valid = PE_118_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_57_io_to_pes_8_out_bits = PE_118_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_57_io_to_pes_9_out_valid = PE_119_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_57_io_to_pes_9_out_bits = PE_119_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_57_io_to_pes_10_out_valid = PE_120_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_57_io_to_pes_10_out_bits = PE_120_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_57_io_to_pes_11_out_valid = PE_121_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_57_io_to_pes_11_out_bits = PE_121_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_57_io_to_pes_12_out_valid = PE_122_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_57_io_to_pes_12_out_bits = PE_122_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_57_io_to_pes_13_out_valid = PE_123_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_57_io_to_pes_13_out_bits = PE_123_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_57_io_to_pes_14_out_valid = PE_124_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_57_io_to_pes_14_out_bits = PE_124_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_57_io_to_pes_15_out_valid = PE_125_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_57_io_to_pes_15_out_bits = PE_125_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_57_io_to_pes_16_out_valid = PE_126_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_57_io_to_pes_16_out_bits = PE_126_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_57_io_to_pes_17_out_valid = PE_127_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_57_io_to_pes_17_out_bits = PE_127_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_57_io_to_pes_18_out_valid = PE_128_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_57_io_to_pes_18_out_bits = PE_128_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_57_io_to_pes_19_out_valid = PE_129_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_57_io_to_pes_19_out_bits = PE_129_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_57_io_to_pes_20_out_valid = PE_130_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_57_io_to_pes_20_out_bits = PE_130_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_57_io_to_pes_21_out_valid = PE_131_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_57_io_to_pes_21_out_bits = PE_131_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_57_io_sig_stat2trans = MultiDimTime_io_index_1 == 16'h0; // @[pe.scala 278:43]
  assign PENetwork_58_clock = clock;
  assign PENetwork_58_reset = reset;
  assign PENetwork_58_io_to_pes_0_out_valid = PE_132_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_58_io_to_pes_0_out_bits = PE_132_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_58_io_to_pes_1_out_valid = PE_133_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_58_io_to_pes_1_out_bits = PE_133_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_58_io_to_pes_2_out_valid = PE_134_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_58_io_to_pes_2_out_bits = PE_134_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_58_io_to_pes_3_out_valid = PE_135_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_58_io_to_pes_3_out_bits = PE_135_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_58_io_to_pes_4_out_valid = PE_136_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_58_io_to_pes_4_out_bits = PE_136_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_58_io_to_pes_5_out_valid = PE_137_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_58_io_to_pes_5_out_bits = PE_137_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_58_io_to_pes_6_out_valid = PE_138_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_58_io_to_pes_6_out_bits = PE_138_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_58_io_to_pes_7_out_valid = PE_139_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_58_io_to_pes_7_out_bits = PE_139_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_58_io_to_pes_8_out_valid = PE_140_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_58_io_to_pes_8_out_bits = PE_140_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_58_io_to_pes_9_out_valid = PE_141_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_58_io_to_pes_9_out_bits = PE_141_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_58_io_to_pes_10_out_valid = PE_142_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_58_io_to_pes_10_out_bits = PE_142_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_58_io_to_pes_11_out_valid = PE_143_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_58_io_to_pes_11_out_bits = PE_143_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_58_io_to_pes_12_out_valid = PE_144_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_58_io_to_pes_12_out_bits = PE_144_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_58_io_to_pes_13_out_valid = PE_145_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_58_io_to_pes_13_out_bits = PE_145_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_58_io_to_pes_14_out_valid = PE_146_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_58_io_to_pes_14_out_bits = PE_146_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_58_io_to_pes_15_out_valid = PE_147_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_58_io_to_pes_15_out_bits = PE_147_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_58_io_to_pes_16_out_valid = PE_148_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_58_io_to_pes_16_out_bits = PE_148_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_58_io_to_pes_17_out_valid = PE_149_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_58_io_to_pes_17_out_bits = PE_149_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_58_io_to_pes_18_out_valid = PE_150_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_58_io_to_pes_18_out_bits = PE_150_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_58_io_to_pes_19_out_valid = PE_151_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_58_io_to_pes_19_out_bits = PE_151_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_58_io_to_pes_20_out_valid = PE_152_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_58_io_to_pes_20_out_bits = PE_152_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_58_io_to_pes_21_out_valid = PE_153_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_58_io_to_pes_21_out_bits = PE_153_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_58_io_sig_stat2trans = MultiDimTime_io_index_1 == 16'h0; // @[pe.scala 278:43]
  assign PENetwork_59_clock = clock;
  assign PENetwork_59_reset = reset;
  assign PENetwork_59_io_to_pes_0_out_valid = PE_154_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_59_io_to_pes_0_out_bits = PE_154_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_59_io_to_pes_1_out_valid = PE_155_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_59_io_to_pes_1_out_bits = PE_155_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_59_io_to_pes_2_out_valid = PE_156_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_59_io_to_pes_2_out_bits = PE_156_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_59_io_to_pes_3_out_valid = PE_157_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_59_io_to_pes_3_out_bits = PE_157_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_59_io_to_pes_4_out_valid = PE_158_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_59_io_to_pes_4_out_bits = PE_158_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_59_io_to_pes_5_out_valid = PE_159_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_59_io_to_pes_5_out_bits = PE_159_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_59_io_to_pes_6_out_valid = PE_160_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_59_io_to_pes_6_out_bits = PE_160_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_59_io_to_pes_7_out_valid = PE_161_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_59_io_to_pes_7_out_bits = PE_161_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_59_io_to_pes_8_out_valid = PE_162_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_59_io_to_pes_8_out_bits = PE_162_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_59_io_to_pes_9_out_valid = PE_163_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_59_io_to_pes_9_out_bits = PE_163_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_59_io_to_pes_10_out_valid = PE_164_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_59_io_to_pes_10_out_bits = PE_164_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_59_io_to_pes_11_out_valid = PE_165_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_59_io_to_pes_11_out_bits = PE_165_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_59_io_to_pes_12_out_valid = PE_166_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_59_io_to_pes_12_out_bits = PE_166_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_59_io_to_pes_13_out_valid = PE_167_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_59_io_to_pes_13_out_bits = PE_167_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_59_io_to_pes_14_out_valid = PE_168_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_59_io_to_pes_14_out_bits = PE_168_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_59_io_to_pes_15_out_valid = PE_169_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_59_io_to_pes_15_out_bits = PE_169_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_59_io_to_pes_16_out_valid = PE_170_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_59_io_to_pes_16_out_bits = PE_170_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_59_io_to_pes_17_out_valid = PE_171_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_59_io_to_pes_17_out_bits = PE_171_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_59_io_to_pes_18_out_valid = PE_172_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_59_io_to_pes_18_out_bits = PE_172_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_59_io_to_pes_19_out_valid = PE_173_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_59_io_to_pes_19_out_bits = PE_173_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_59_io_to_pes_20_out_valid = PE_174_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_59_io_to_pes_20_out_bits = PE_174_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_59_io_to_pes_21_out_valid = PE_175_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_59_io_to_pes_21_out_bits = PE_175_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_59_io_sig_stat2trans = MultiDimTime_io_index_1 == 16'h0; // @[pe.scala 278:43]
  assign PENetwork_60_clock = clock;
  assign PENetwork_60_reset = reset;
  assign PENetwork_60_io_to_pes_0_out_valid = PE_176_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_60_io_to_pes_0_out_bits = PE_176_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_60_io_to_pes_1_out_valid = PE_177_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_60_io_to_pes_1_out_bits = PE_177_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_60_io_to_pes_2_out_valid = PE_178_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_60_io_to_pes_2_out_bits = PE_178_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_60_io_to_pes_3_out_valid = PE_179_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_60_io_to_pes_3_out_bits = PE_179_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_60_io_to_pes_4_out_valid = PE_180_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_60_io_to_pes_4_out_bits = PE_180_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_60_io_to_pes_5_out_valid = PE_181_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_60_io_to_pes_5_out_bits = PE_181_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_60_io_to_pes_6_out_valid = PE_182_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_60_io_to_pes_6_out_bits = PE_182_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_60_io_to_pes_7_out_valid = PE_183_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_60_io_to_pes_7_out_bits = PE_183_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_60_io_to_pes_8_out_valid = PE_184_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_60_io_to_pes_8_out_bits = PE_184_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_60_io_to_pes_9_out_valid = PE_185_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_60_io_to_pes_9_out_bits = PE_185_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_60_io_to_pes_10_out_valid = PE_186_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_60_io_to_pes_10_out_bits = PE_186_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_60_io_to_pes_11_out_valid = PE_187_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_60_io_to_pes_11_out_bits = PE_187_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_60_io_to_pes_12_out_valid = PE_188_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_60_io_to_pes_12_out_bits = PE_188_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_60_io_to_pes_13_out_valid = PE_189_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_60_io_to_pes_13_out_bits = PE_189_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_60_io_to_pes_14_out_valid = PE_190_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_60_io_to_pes_14_out_bits = PE_190_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_60_io_to_pes_15_out_valid = PE_191_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_60_io_to_pes_15_out_bits = PE_191_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_60_io_to_pes_16_out_valid = PE_192_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_60_io_to_pes_16_out_bits = PE_192_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_60_io_to_pes_17_out_valid = PE_193_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_60_io_to_pes_17_out_bits = PE_193_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_60_io_to_pes_18_out_valid = PE_194_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_60_io_to_pes_18_out_bits = PE_194_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_60_io_to_pes_19_out_valid = PE_195_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_60_io_to_pes_19_out_bits = PE_195_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_60_io_to_pes_20_out_valid = PE_196_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_60_io_to_pes_20_out_bits = PE_196_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_60_io_to_pes_21_out_valid = PE_197_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_60_io_to_pes_21_out_bits = PE_197_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_60_io_sig_stat2trans = MultiDimTime_io_index_1 == 16'h0; // @[pe.scala 278:43]
  assign PENetwork_61_clock = clock;
  assign PENetwork_61_reset = reset;
  assign PENetwork_61_io_to_pes_0_out_valid = PE_198_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_61_io_to_pes_0_out_bits = PE_198_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_61_io_to_pes_1_out_valid = PE_199_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_61_io_to_pes_1_out_bits = PE_199_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_61_io_to_pes_2_out_valid = PE_200_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_61_io_to_pes_2_out_bits = PE_200_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_61_io_to_pes_3_out_valid = PE_201_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_61_io_to_pes_3_out_bits = PE_201_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_61_io_to_pes_4_out_valid = PE_202_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_61_io_to_pes_4_out_bits = PE_202_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_61_io_to_pes_5_out_valid = PE_203_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_61_io_to_pes_5_out_bits = PE_203_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_61_io_to_pes_6_out_valid = PE_204_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_61_io_to_pes_6_out_bits = PE_204_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_61_io_to_pes_7_out_valid = PE_205_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_61_io_to_pes_7_out_bits = PE_205_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_61_io_to_pes_8_out_valid = PE_206_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_61_io_to_pes_8_out_bits = PE_206_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_61_io_to_pes_9_out_valid = PE_207_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_61_io_to_pes_9_out_bits = PE_207_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_61_io_to_pes_10_out_valid = PE_208_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_61_io_to_pes_10_out_bits = PE_208_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_61_io_to_pes_11_out_valid = PE_209_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_61_io_to_pes_11_out_bits = PE_209_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_61_io_to_pes_12_out_valid = PE_210_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_61_io_to_pes_12_out_bits = PE_210_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_61_io_to_pes_13_out_valid = PE_211_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_61_io_to_pes_13_out_bits = PE_211_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_61_io_to_pes_14_out_valid = PE_212_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_61_io_to_pes_14_out_bits = PE_212_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_61_io_to_pes_15_out_valid = PE_213_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_61_io_to_pes_15_out_bits = PE_213_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_61_io_to_pes_16_out_valid = PE_214_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_61_io_to_pes_16_out_bits = PE_214_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_61_io_to_pes_17_out_valid = PE_215_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_61_io_to_pes_17_out_bits = PE_215_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_61_io_to_pes_18_out_valid = PE_216_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_61_io_to_pes_18_out_bits = PE_216_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_61_io_to_pes_19_out_valid = PE_217_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_61_io_to_pes_19_out_bits = PE_217_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_61_io_to_pes_20_out_valid = PE_218_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_61_io_to_pes_20_out_bits = PE_218_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_61_io_to_pes_21_out_valid = PE_219_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_61_io_to_pes_21_out_bits = PE_219_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_61_io_sig_stat2trans = MultiDimTime_io_index_1 == 16'h0; // @[pe.scala 278:43]
  assign PENetwork_62_clock = clock;
  assign PENetwork_62_reset = reset;
  assign PENetwork_62_io_to_pes_0_out_valid = PE_220_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_62_io_to_pes_0_out_bits = PE_220_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_62_io_to_pes_1_out_valid = PE_221_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_62_io_to_pes_1_out_bits = PE_221_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_62_io_to_pes_2_out_valid = PE_222_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_62_io_to_pes_2_out_bits = PE_222_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_62_io_to_pes_3_out_valid = PE_223_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_62_io_to_pes_3_out_bits = PE_223_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_62_io_to_pes_4_out_valid = PE_224_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_62_io_to_pes_4_out_bits = PE_224_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_62_io_to_pes_5_out_valid = PE_225_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_62_io_to_pes_5_out_bits = PE_225_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_62_io_to_pes_6_out_valid = PE_226_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_62_io_to_pes_6_out_bits = PE_226_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_62_io_to_pes_7_out_valid = PE_227_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_62_io_to_pes_7_out_bits = PE_227_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_62_io_to_pes_8_out_valid = PE_228_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_62_io_to_pes_8_out_bits = PE_228_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_62_io_to_pes_9_out_valid = PE_229_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_62_io_to_pes_9_out_bits = PE_229_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_62_io_to_pes_10_out_valid = PE_230_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_62_io_to_pes_10_out_bits = PE_230_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_62_io_to_pes_11_out_valid = PE_231_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_62_io_to_pes_11_out_bits = PE_231_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_62_io_to_pes_12_out_valid = PE_232_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_62_io_to_pes_12_out_bits = PE_232_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_62_io_to_pes_13_out_valid = PE_233_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_62_io_to_pes_13_out_bits = PE_233_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_62_io_to_pes_14_out_valid = PE_234_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_62_io_to_pes_14_out_bits = PE_234_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_62_io_to_pes_15_out_valid = PE_235_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_62_io_to_pes_15_out_bits = PE_235_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_62_io_to_pes_16_out_valid = PE_236_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_62_io_to_pes_16_out_bits = PE_236_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_62_io_to_pes_17_out_valid = PE_237_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_62_io_to_pes_17_out_bits = PE_237_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_62_io_to_pes_18_out_valid = PE_238_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_62_io_to_pes_18_out_bits = PE_238_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_62_io_to_pes_19_out_valid = PE_239_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_62_io_to_pes_19_out_bits = PE_239_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_62_io_to_pes_20_out_valid = PE_240_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_62_io_to_pes_20_out_bits = PE_240_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_62_io_to_pes_21_out_valid = PE_241_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_62_io_to_pes_21_out_bits = PE_241_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_62_io_sig_stat2trans = MultiDimTime_io_index_1 == 16'h0; // @[pe.scala 278:43]
  assign PENetwork_63_clock = clock;
  assign PENetwork_63_reset = reset;
  assign PENetwork_63_io_to_pes_0_out_valid = PE_242_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_63_io_to_pes_0_out_bits = PE_242_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_63_io_to_pes_1_out_valid = PE_243_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_63_io_to_pes_1_out_bits = PE_243_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_63_io_to_pes_2_out_valid = PE_244_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_63_io_to_pes_2_out_bits = PE_244_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_63_io_to_pes_3_out_valid = PE_245_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_63_io_to_pes_3_out_bits = PE_245_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_63_io_to_pes_4_out_valid = PE_246_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_63_io_to_pes_4_out_bits = PE_246_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_63_io_to_pes_5_out_valid = PE_247_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_63_io_to_pes_5_out_bits = PE_247_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_63_io_to_pes_6_out_valid = PE_248_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_63_io_to_pes_6_out_bits = PE_248_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_63_io_to_pes_7_out_valid = PE_249_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_63_io_to_pes_7_out_bits = PE_249_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_63_io_to_pes_8_out_valid = PE_250_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_63_io_to_pes_8_out_bits = PE_250_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_63_io_to_pes_9_out_valid = PE_251_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_63_io_to_pes_9_out_bits = PE_251_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_63_io_to_pes_10_out_valid = PE_252_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_63_io_to_pes_10_out_bits = PE_252_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_63_io_to_pes_11_out_valid = PE_253_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_63_io_to_pes_11_out_bits = PE_253_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_63_io_to_pes_12_out_valid = PE_254_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_63_io_to_pes_12_out_bits = PE_254_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_63_io_to_pes_13_out_valid = PE_255_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_63_io_to_pes_13_out_bits = PE_255_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_63_io_to_pes_14_out_valid = PE_256_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_63_io_to_pes_14_out_bits = PE_256_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_63_io_to_pes_15_out_valid = PE_257_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_63_io_to_pes_15_out_bits = PE_257_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_63_io_to_pes_16_out_valid = PE_258_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_63_io_to_pes_16_out_bits = PE_258_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_63_io_to_pes_17_out_valid = PE_259_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_63_io_to_pes_17_out_bits = PE_259_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_63_io_to_pes_18_out_valid = PE_260_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_63_io_to_pes_18_out_bits = PE_260_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_63_io_to_pes_19_out_valid = PE_261_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_63_io_to_pes_19_out_bits = PE_261_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_63_io_to_pes_20_out_valid = PE_262_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_63_io_to_pes_20_out_bits = PE_262_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_63_io_to_pes_21_out_valid = PE_263_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_63_io_to_pes_21_out_bits = PE_263_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_63_io_sig_stat2trans = MultiDimTime_io_index_1 == 16'h0; // @[pe.scala 278:43]
  assign PENetwork_64_clock = clock;
  assign PENetwork_64_reset = reset;
  assign PENetwork_64_io_to_pes_0_out_valid = PE_264_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_64_io_to_pes_0_out_bits = PE_264_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_64_io_to_pes_1_out_valid = PE_265_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_64_io_to_pes_1_out_bits = PE_265_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_64_io_to_pes_2_out_valid = PE_266_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_64_io_to_pes_2_out_bits = PE_266_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_64_io_to_pes_3_out_valid = PE_267_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_64_io_to_pes_3_out_bits = PE_267_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_64_io_to_pes_4_out_valid = PE_268_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_64_io_to_pes_4_out_bits = PE_268_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_64_io_to_pes_5_out_valid = PE_269_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_64_io_to_pes_5_out_bits = PE_269_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_64_io_to_pes_6_out_valid = PE_270_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_64_io_to_pes_6_out_bits = PE_270_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_64_io_to_pes_7_out_valid = PE_271_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_64_io_to_pes_7_out_bits = PE_271_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_64_io_to_pes_8_out_valid = PE_272_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_64_io_to_pes_8_out_bits = PE_272_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_64_io_to_pes_9_out_valid = PE_273_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_64_io_to_pes_9_out_bits = PE_273_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_64_io_to_pes_10_out_valid = PE_274_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_64_io_to_pes_10_out_bits = PE_274_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_64_io_to_pes_11_out_valid = PE_275_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_64_io_to_pes_11_out_bits = PE_275_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_64_io_to_pes_12_out_valid = PE_276_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_64_io_to_pes_12_out_bits = PE_276_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_64_io_to_pes_13_out_valid = PE_277_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_64_io_to_pes_13_out_bits = PE_277_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_64_io_to_pes_14_out_valid = PE_278_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_64_io_to_pes_14_out_bits = PE_278_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_64_io_to_pes_15_out_valid = PE_279_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_64_io_to_pes_15_out_bits = PE_279_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_64_io_to_pes_16_out_valid = PE_280_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_64_io_to_pes_16_out_bits = PE_280_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_64_io_to_pes_17_out_valid = PE_281_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_64_io_to_pes_17_out_bits = PE_281_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_64_io_to_pes_18_out_valid = PE_282_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_64_io_to_pes_18_out_bits = PE_282_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_64_io_to_pes_19_out_valid = PE_283_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_64_io_to_pes_19_out_bits = PE_283_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_64_io_to_pes_20_out_valid = PE_284_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_64_io_to_pes_20_out_bits = PE_284_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_64_io_to_pes_21_out_valid = PE_285_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_64_io_to_pes_21_out_bits = PE_285_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_64_io_sig_stat2trans = MultiDimTime_io_index_1 == 16'h0; // @[pe.scala 278:43]
  assign PENetwork_65_clock = clock;
  assign PENetwork_65_reset = reset;
  assign PENetwork_65_io_to_pes_0_out_valid = PE_286_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_65_io_to_pes_0_out_bits = PE_286_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_65_io_to_pes_1_out_valid = PE_287_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_65_io_to_pes_1_out_bits = PE_287_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_65_io_to_pes_2_out_valid = PE_288_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_65_io_to_pes_2_out_bits = PE_288_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_65_io_to_pes_3_out_valid = PE_289_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_65_io_to_pes_3_out_bits = PE_289_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_65_io_to_pes_4_out_valid = PE_290_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_65_io_to_pes_4_out_bits = PE_290_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_65_io_to_pes_5_out_valid = PE_291_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_65_io_to_pes_5_out_bits = PE_291_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_65_io_to_pes_6_out_valid = PE_292_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_65_io_to_pes_6_out_bits = PE_292_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_65_io_to_pes_7_out_valid = PE_293_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_65_io_to_pes_7_out_bits = PE_293_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_65_io_to_pes_8_out_valid = PE_294_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_65_io_to_pes_8_out_bits = PE_294_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_65_io_to_pes_9_out_valid = PE_295_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_65_io_to_pes_9_out_bits = PE_295_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_65_io_to_pes_10_out_valid = PE_296_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_65_io_to_pes_10_out_bits = PE_296_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_65_io_to_pes_11_out_valid = PE_297_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_65_io_to_pes_11_out_bits = PE_297_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_65_io_to_pes_12_out_valid = PE_298_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_65_io_to_pes_12_out_bits = PE_298_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_65_io_to_pes_13_out_valid = PE_299_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_65_io_to_pes_13_out_bits = PE_299_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_65_io_to_pes_14_out_valid = PE_300_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_65_io_to_pes_14_out_bits = PE_300_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_65_io_to_pes_15_out_valid = PE_301_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_65_io_to_pes_15_out_bits = PE_301_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_65_io_to_pes_16_out_valid = PE_302_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_65_io_to_pes_16_out_bits = PE_302_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_65_io_to_pes_17_out_valid = PE_303_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_65_io_to_pes_17_out_bits = PE_303_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_65_io_to_pes_18_out_valid = PE_304_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_65_io_to_pes_18_out_bits = PE_304_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_65_io_to_pes_19_out_valid = PE_305_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_65_io_to_pes_19_out_bits = PE_305_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_65_io_to_pes_20_out_valid = PE_306_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_65_io_to_pes_20_out_bits = PE_306_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_65_io_to_pes_21_out_valid = PE_307_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_65_io_to_pes_21_out_bits = PE_307_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_65_io_sig_stat2trans = MultiDimTime_io_index_1 == 16'h0; // @[pe.scala 278:43]
  assign PENetwork_66_clock = clock;
  assign PENetwork_66_reset = reset;
  assign PENetwork_66_io_to_pes_0_out_valid = PE_308_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_66_io_to_pes_0_out_bits = PE_308_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_66_io_to_pes_1_out_valid = PE_309_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_66_io_to_pes_1_out_bits = PE_309_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_66_io_to_pes_2_out_valid = PE_310_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_66_io_to_pes_2_out_bits = PE_310_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_66_io_to_pes_3_out_valid = PE_311_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_66_io_to_pes_3_out_bits = PE_311_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_66_io_to_pes_4_out_valid = PE_312_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_66_io_to_pes_4_out_bits = PE_312_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_66_io_to_pes_5_out_valid = PE_313_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_66_io_to_pes_5_out_bits = PE_313_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_66_io_to_pes_6_out_valid = PE_314_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_66_io_to_pes_6_out_bits = PE_314_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_66_io_to_pes_7_out_valid = PE_315_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_66_io_to_pes_7_out_bits = PE_315_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_66_io_to_pes_8_out_valid = PE_316_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_66_io_to_pes_8_out_bits = PE_316_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_66_io_to_pes_9_out_valid = PE_317_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_66_io_to_pes_9_out_bits = PE_317_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_66_io_to_pes_10_out_valid = PE_318_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_66_io_to_pes_10_out_bits = PE_318_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_66_io_to_pes_11_out_valid = PE_319_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_66_io_to_pes_11_out_bits = PE_319_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_66_io_to_pes_12_out_valid = PE_320_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_66_io_to_pes_12_out_bits = PE_320_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_66_io_to_pes_13_out_valid = PE_321_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_66_io_to_pes_13_out_bits = PE_321_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_66_io_to_pes_14_out_valid = PE_322_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_66_io_to_pes_14_out_bits = PE_322_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_66_io_to_pes_15_out_valid = PE_323_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_66_io_to_pes_15_out_bits = PE_323_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_66_io_to_pes_16_out_valid = PE_324_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_66_io_to_pes_16_out_bits = PE_324_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_66_io_to_pes_17_out_valid = PE_325_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_66_io_to_pes_17_out_bits = PE_325_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_66_io_to_pes_18_out_valid = PE_326_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_66_io_to_pes_18_out_bits = PE_326_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_66_io_to_pes_19_out_valid = PE_327_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_66_io_to_pes_19_out_bits = PE_327_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_66_io_to_pes_20_out_valid = PE_328_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_66_io_to_pes_20_out_bits = PE_328_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_66_io_to_pes_21_out_valid = PE_329_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_66_io_to_pes_21_out_bits = PE_329_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_66_io_sig_stat2trans = MultiDimTime_io_index_1 == 16'h0; // @[pe.scala 278:43]
  assign PENetwork_67_clock = clock;
  assign PENetwork_67_reset = reset;
  assign PENetwork_67_io_to_pes_0_out_valid = PE_330_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_67_io_to_pes_0_out_bits = PE_330_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_67_io_to_pes_1_out_valid = PE_331_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_67_io_to_pes_1_out_bits = PE_331_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_67_io_to_pes_2_out_valid = PE_332_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_67_io_to_pes_2_out_bits = PE_332_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_67_io_to_pes_3_out_valid = PE_333_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_67_io_to_pes_3_out_bits = PE_333_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_67_io_to_pes_4_out_valid = PE_334_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_67_io_to_pes_4_out_bits = PE_334_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_67_io_to_pes_5_out_valid = PE_335_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_67_io_to_pes_5_out_bits = PE_335_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_67_io_to_pes_6_out_valid = PE_336_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_67_io_to_pes_6_out_bits = PE_336_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_67_io_to_pes_7_out_valid = PE_337_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_67_io_to_pes_7_out_bits = PE_337_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_67_io_to_pes_8_out_valid = PE_338_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_67_io_to_pes_8_out_bits = PE_338_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_67_io_to_pes_9_out_valid = PE_339_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_67_io_to_pes_9_out_bits = PE_339_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_67_io_to_pes_10_out_valid = PE_340_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_67_io_to_pes_10_out_bits = PE_340_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_67_io_to_pes_11_out_valid = PE_341_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_67_io_to_pes_11_out_bits = PE_341_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_67_io_to_pes_12_out_valid = PE_342_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_67_io_to_pes_12_out_bits = PE_342_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_67_io_to_pes_13_out_valid = PE_343_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_67_io_to_pes_13_out_bits = PE_343_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_67_io_to_pes_14_out_valid = PE_344_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_67_io_to_pes_14_out_bits = PE_344_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_67_io_to_pes_15_out_valid = PE_345_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_67_io_to_pes_15_out_bits = PE_345_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_67_io_to_pes_16_out_valid = PE_346_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_67_io_to_pes_16_out_bits = PE_346_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_67_io_to_pes_17_out_valid = PE_347_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_67_io_to_pes_17_out_bits = PE_347_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_67_io_to_pes_18_out_valid = PE_348_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_67_io_to_pes_18_out_bits = PE_348_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_67_io_to_pes_19_out_valid = PE_349_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_67_io_to_pes_19_out_bits = PE_349_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_67_io_to_pes_20_out_valid = PE_350_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_67_io_to_pes_20_out_bits = PE_350_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_67_io_to_pes_21_out_valid = PE_351_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_67_io_to_pes_21_out_bits = PE_351_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_67_io_sig_stat2trans = MultiDimTime_io_index_1 == 16'h0; // @[pe.scala 278:43]
  assign PENetwork_68_clock = clock;
  assign PENetwork_68_reset = reset;
  assign PENetwork_68_io_to_pes_0_out_valid = PE_352_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_68_io_to_pes_0_out_bits = PE_352_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_68_io_to_pes_1_out_valid = PE_353_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_68_io_to_pes_1_out_bits = PE_353_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_68_io_to_pes_2_out_valid = PE_354_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_68_io_to_pes_2_out_bits = PE_354_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_68_io_to_pes_3_out_valid = PE_355_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_68_io_to_pes_3_out_bits = PE_355_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_68_io_to_pes_4_out_valid = PE_356_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_68_io_to_pes_4_out_bits = PE_356_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_68_io_to_pes_5_out_valid = PE_357_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_68_io_to_pes_5_out_bits = PE_357_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_68_io_to_pes_6_out_valid = PE_358_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_68_io_to_pes_6_out_bits = PE_358_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_68_io_to_pes_7_out_valid = PE_359_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_68_io_to_pes_7_out_bits = PE_359_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_68_io_to_pes_8_out_valid = PE_360_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_68_io_to_pes_8_out_bits = PE_360_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_68_io_to_pes_9_out_valid = PE_361_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_68_io_to_pes_9_out_bits = PE_361_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_68_io_to_pes_10_out_valid = PE_362_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_68_io_to_pes_10_out_bits = PE_362_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_68_io_to_pes_11_out_valid = PE_363_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_68_io_to_pes_11_out_bits = PE_363_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_68_io_to_pes_12_out_valid = PE_364_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_68_io_to_pes_12_out_bits = PE_364_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_68_io_to_pes_13_out_valid = PE_365_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_68_io_to_pes_13_out_bits = PE_365_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_68_io_to_pes_14_out_valid = PE_366_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_68_io_to_pes_14_out_bits = PE_366_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_68_io_to_pes_15_out_valid = PE_367_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_68_io_to_pes_15_out_bits = PE_367_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_68_io_to_pes_16_out_valid = PE_368_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_68_io_to_pes_16_out_bits = PE_368_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_68_io_to_pes_17_out_valid = PE_369_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_68_io_to_pes_17_out_bits = PE_369_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_68_io_to_pes_18_out_valid = PE_370_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_68_io_to_pes_18_out_bits = PE_370_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_68_io_to_pes_19_out_valid = PE_371_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_68_io_to_pes_19_out_bits = PE_371_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_68_io_to_pes_20_out_valid = PE_372_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_68_io_to_pes_20_out_bits = PE_372_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_68_io_to_pes_21_out_valid = PE_373_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_68_io_to_pes_21_out_bits = PE_373_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_68_io_sig_stat2trans = MultiDimTime_io_index_1 == 16'h0; // @[pe.scala 278:43]
  assign PENetwork_69_clock = clock;
  assign PENetwork_69_reset = reset;
  assign PENetwork_69_io_to_pes_0_out_valid = PE_374_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_69_io_to_pes_0_out_bits = PE_374_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_69_io_to_pes_1_out_valid = PE_375_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_69_io_to_pes_1_out_bits = PE_375_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_69_io_to_pes_2_out_valid = PE_376_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_69_io_to_pes_2_out_bits = PE_376_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_69_io_to_pes_3_out_valid = PE_377_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_69_io_to_pes_3_out_bits = PE_377_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_69_io_to_pes_4_out_valid = PE_378_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_69_io_to_pes_4_out_bits = PE_378_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_69_io_to_pes_5_out_valid = PE_379_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_69_io_to_pes_5_out_bits = PE_379_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_69_io_to_pes_6_out_valid = PE_380_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_69_io_to_pes_6_out_bits = PE_380_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_69_io_to_pes_7_out_valid = PE_381_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_69_io_to_pes_7_out_bits = PE_381_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_69_io_to_pes_8_out_valid = PE_382_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_69_io_to_pes_8_out_bits = PE_382_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_69_io_to_pes_9_out_valid = PE_383_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_69_io_to_pes_9_out_bits = PE_383_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_69_io_to_pes_10_out_valid = PE_384_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_69_io_to_pes_10_out_bits = PE_384_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_69_io_to_pes_11_out_valid = PE_385_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_69_io_to_pes_11_out_bits = PE_385_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_69_io_to_pes_12_out_valid = PE_386_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_69_io_to_pes_12_out_bits = PE_386_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_69_io_to_pes_13_out_valid = PE_387_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_69_io_to_pes_13_out_bits = PE_387_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_69_io_to_pes_14_out_valid = PE_388_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_69_io_to_pes_14_out_bits = PE_388_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_69_io_to_pes_15_out_valid = PE_389_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_69_io_to_pes_15_out_bits = PE_389_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_69_io_to_pes_16_out_valid = PE_390_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_69_io_to_pes_16_out_bits = PE_390_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_69_io_to_pes_17_out_valid = PE_391_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_69_io_to_pes_17_out_bits = PE_391_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_69_io_to_pes_18_out_valid = PE_392_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_69_io_to_pes_18_out_bits = PE_392_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_69_io_to_pes_19_out_valid = PE_393_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_69_io_to_pes_19_out_bits = PE_393_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_69_io_to_pes_20_out_valid = PE_394_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_69_io_to_pes_20_out_bits = PE_394_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_69_io_to_pes_21_out_valid = PE_395_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_69_io_to_pes_21_out_bits = PE_395_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_69_io_sig_stat2trans = MultiDimTime_io_index_1 == 16'h0; // @[pe.scala 278:43]
  assign PENetwork_70_clock = clock;
  assign PENetwork_70_reset = reset;
  assign PENetwork_70_io_to_pes_0_out_valid = PE_396_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_70_io_to_pes_0_out_bits = PE_396_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_70_io_to_pes_1_out_valid = PE_397_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_70_io_to_pes_1_out_bits = PE_397_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_70_io_to_pes_2_out_valid = PE_398_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_70_io_to_pes_2_out_bits = PE_398_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_70_io_to_pes_3_out_valid = PE_399_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_70_io_to_pes_3_out_bits = PE_399_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_70_io_to_pes_4_out_valid = PE_400_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_70_io_to_pes_4_out_bits = PE_400_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_70_io_to_pes_5_out_valid = PE_401_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_70_io_to_pes_5_out_bits = PE_401_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_70_io_to_pes_6_out_valid = PE_402_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_70_io_to_pes_6_out_bits = PE_402_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_70_io_to_pes_7_out_valid = PE_403_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_70_io_to_pes_7_out_bits = PE_403_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_70_io_to_pes_8_out_valid = PE_404_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_70_io_to_pes_8_out_bits = PE_404_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_70_io_to_pes_9_out_valid = PE_405_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_70_io_to_pes_9_out_bits = PE_405_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_70_io_to_pes_10_out_valid = PE_406_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_70_io_to_pes_10_out_bits = PE_406_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_70_io_to_pes_11_out_valid = PE_407_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_70_io_to_pes_11_out_bits = PE_407_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_70_io_to_pes_12_out_valid = PE_408_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_70_io_to_pes_12_out_bits = PE_408_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_70_io_to_pes_13_out_valid = PE_409_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_70_io_to_pes_13_out_bits = PE_409_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_70_io_to_pes_14_out_valid = PE_410_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_70_io_to_pes_14_out_bits = PE_410_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_70_io_to_pes_15_out_valid = PE_411_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_70_io_to_pes_15_out_bits = PE_411_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_70_io_to_pes_16_out_valid = PE_412_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_70_io_to_pes_16_out_bits = PE_412_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_70_io_to_pes_17_out_valid = PE_413_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_70_io_to_pes_17_out_bits = PE_413_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_70_io_to_pes_18_out_valid = PE_414_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_70_io_to_pes_18_out_bits = PE_414_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_70_io_to_pes_19_out_valid = PE_415_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_70_io_to_pes_19_out_bits = PE_415_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_70_io_to_pes_20_out_valid = PE_416_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_70_io_to_pes_20_out_bits = PE_416_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_70_io_to_pes_21_out_valid = PE_417_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_70_io_to_pes_21_out_bits = PE_417_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_70_io_sig_stat2trans = MultiDimTime_io_index_1 == 16'h0; // @[pe.scala 278:43]
  assign PENetwork_71_clock = clock;
  assign PENetwork_71_reset = reset;
  assign PENetwork_71_io_to_pes_0_out_valid = PE_418_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_71_io_to_pes_0_out_bits = PE_418_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_71_io_to_pes_1_out_valid = PE_419_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_71_io_to_pes_1_out_bits = PE_419_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_71_io_to_pes_2_out_valid = PE_420_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_71_io_to_pes_2_out_bits = PE_420_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_71_io_to_pes_3_out_valid = PE_421_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_71_io_to_pes_3_out_bits = PE_421_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_71_io_to_pes_4_out_valid = PE_422_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_71_io_to_pes_4_out_bits = PE_422_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_71_io_to_pes_5_out_valid = PE_423_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_71_io_to_pes_5_out_bits = PE_423_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_71_io_to_pes_6_out_valid = PE_424_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_71_io_to_pes_6_out_bits = PE_424_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_71_io_to_pes_7_out_valid = PE_425_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_71_io_to_pes_7_out_bits = PE_425_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_71_io_to_pes_8_out_valid = PE_426_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_71_io_to_pes_8_out_bits = PE_426_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_71_io_to_pes_9_out_valid = PE_427_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_71_io_to_pes_9_out_bits = PE_427_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_71_io_to_pes_10_out_valid = PE_428_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_71_io_to_pes_10_out_bits = PE_428_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_71_io_to_pes_11_out_valid = PE_429_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_71_io_to_pes_11_out_bits = PE_429_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_71_io_to_pes_12_out_valid = PE_430_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_71_io_to_pes_12_out_bits = PE_430_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_71_io_to_pes_13_out_valid = PE_431_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_71_io_to_pes_13_out_bits = PE_431_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_71_io_to_pes_14_out_valid = PE_432_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_71_io_to_pes_14_out_bits = PE_432_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_71_io_to_pes_15_out_valid = PE_433_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_71_io_to_pes_15_out_bits = PE_433_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_71_io_to_pes_16_out_valid = PE_434_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_71_io_to_pes_16_out_bits = PE_434_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_71_io_to_pes_17_out_valid = PE_435_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_71_io_to_pes_17_out_bits = PE_435_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_71_io_to_pes_18_out_valid = PE_436_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_71_io_to_pes_18_out_bits = PE_436_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_71_io_to_pes_19_out_valid = PE_437_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_71_io_to_pes_19_out_bits = PE_437_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_71_io_to_pes_20_out_valid = PE_438_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_71_io_to_pes_20_out_bits = PE_438_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_71_io_to_pes_21_out_valid = PE_439_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_71_io_to_pes_21_out_bits = PE_439_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_71_io_sig_stat2trans = MultiDimTime_io_index_1 == 16'h0; // @[pe.scala 278:43]
  assign PENetwork_72_clock = clock;
  assign PENetwork_72_reset = reset;
  assign PENetwork_72_io_to_pes_0_out_valid = PE_440_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_72_io_to_pes_0_out_bits = PE_440_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_72_io_to_pes_1_out_valid = PE_441_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_72_io_to_pes_1_out_bits = PE_441_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_72_io_to_pes_2_out_valid = PE_442_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_72_io_to_pes_2_out_bits = PE_442_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_72_io_to_pes_3_out_valid = PE_443_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_72_io_to_pes_3_out_bits = PE_443_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_72_io_to_pes_4_out_valid = PE_444_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_72_io_to_pes_4_out_bits = PE_444_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_72_io_to_pes_5_out_valid = PE_445_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_72_io_to_pes_5_out_bits = PE_445_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_72_io_to_pes_6_out_valid = PE_446_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_72_io_to_pes_6_out_bits = PE_446_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_72_io_to_pes_7_out_valid = PE_447_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_72_io_to_pes_7_out_bits = PE_447_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_72_io_to_pes_8_out_valid = PE_448_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_72_io_to_pes_8_out_bits = PE_448_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_72_io_to_pes_9_out_valid = PE_449_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_72_io_to_pes_9_out_bits = PE_449_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_72_io_to_pes_10_out_valid = PE_450_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_72_io_to_pes_10_out_bits = PE_450_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_72_io_to_pes_11_out_valid = PE_451_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_72_io_to_pes_11_out_bits = PE_451_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_72_io_to_pes_12_out_valid = PE_452_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_72_io_to_pes_12_out_bits = PE_452_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_72_io_to_pes_13_out_valid = PE_453_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_72_io_to_pes_13_out_bits = PE_453_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_72_io_to_pes_14_out_valid = PE_454_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_72_io_to_pes_14_out_bits = PE_454_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_72_io_to_pes_15_out_valid = PE_455_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_72_io_to_pes_15_out_bits = PE_455_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_72_io_to_pes_16_out_valid = PE_456_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_72_io_to_pes_16_out_bits = PE_456_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_72_io_to_pes_17_out_valid = PE_457_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_72_io_to_pes_17_out_bits = PE_457_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_72_io_to_pes_18_out_valid = PE_458_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_72_io_to_pes_18_out_bits = PE_458_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_72_io_to_pes_19_out_valid = PE_459_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_72_io_to_pes_19_out_bits = PE_459_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_72_io_to_pes_20_out_valid = PE_460_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_72_io_to_pes_20_out_bits = PE_460_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_72_io_to_pes_21_out_valid = PE_461_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_72_io_to_pes_21_out_bits = PE_461_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_72_io_sig_stat2trans = MultiDimTime_io_index_1 == 16'h0; // @[pe.scala 278:43]
  assign PENetwork_73_clock = clock;
  assign PENetwork_73_reset = reset;
  assign PENetwork_73_io_to_pes_0_out_valid = PE_462_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_73_io_to_pes_0_out_bits = PE_462_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_73_io_to_pes_1_out_valid = PE_463_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_73_io_to_pes_1_out_bits = PE_463_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_73_io_to_pes_2_out_valid = PE_464_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_73_io_to_pes_2_out_bits = PE_464_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_73_io_to_pes_3_out_valid = PE_465_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_73_io_to_pes_3_out_bits = PE_465_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_73_io_to_pes_4_out_valid = PE_466_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_73_io_to_pes_4_out_bits = PE_466_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_73_io_to_pes_5_out_valid = PE_467_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_73_io_to_pes_5_out_bits = PE_467_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_73_io_to_pes_6_out_valid = PE_468_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_73_io_to_pes_6_out_bits = PE_468_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_73_io_to_pes_7_out_valid = PE_469_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_73_io_to_pes_7_out_bits = PE_469_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_73_io_to_pes_8_out_valid = PE_470_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_73_io_to_pes_8_out_bits = PE_470_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_73_io_to_pes_9_out_valid = PE_471_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_73_io_to_pes_9_out_bits = PE_471_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_73_io_to_pes_10_out_valid = PE_472_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_73_io_to_pes_10_out_bits = PE_472_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_73_io_to_pes_11_out_valid = PE_473_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_73_io_to_pes_11_out_bits = PE_473_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_73_io_to_pes_12_out_valid = PE_474_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_73_io_to_pes_12_out_bits = PE_474_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_73_io_to_pes_13_out_valid = PE_475_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_73_io_to_pes_13_out_bits = PE_475_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_73_io_to_pes_14_out_valid = PE_476_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_73_io_to_pes_14_out_bits = PE_476_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_73_io_to_pes_15_out_valid = PE_477_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_73_io_to_pes_15_out_bits = PE_477_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_73_io_to_pes_16_out_valid = PE_478_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_73_io_to_pes_16_out_bits = PE_478_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_73_io_to_pes_17_out_valid = PE_479_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_73_io_to_pes_17_out_bits = PE_479_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_73_io_to_pes_18_out_valid = PE_480_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_73_io_to_pes_18_out_bits = PE_480_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_73_io_to_pes_19_out_valid = PE_481_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_73_io_to_pes_19_out_bits = PE_481_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_73_io_to_pes_20_out_valid = PE_482_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_73_io_to_pes_20_out_bits = PE_482_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_73_io_to_pes_21_out_valid = PE_483_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_73_io_to_pes_21_out_bits = PE_483_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_73_io_sig_stat2trans = MultiDimTime_io_index_1 == 16'h0; // @[pe.scala 278:43]
  assign PENetwork_74_clock = clock;
  assign PENetwork_74_reset = reset;
  assign PENetwork_74_io_to_pes_0_out_valid = PE_484_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_74_io_to_pes_0_out_bits = PE_484_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_74_io_to_pes_1_out_valid = PE_485_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_74_io_to_pes_1_out_bits = PE_485_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_74_io_to_pes_2_out_valid = PE_486_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_74_io_to_pes_2_out_bits = PE_486_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_74_io_to_pes_3_out_valid = PE_487_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_74_io_to_pes_3_out_bits = PE_487_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_74_io_to_pes_4_out_valid = PE_488_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_74_io_to_pes_4_out_bits = PE_488_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_74_io_to_pes_5_out_valid = PE_489_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_74_io_to_pes_5_out_bits = PE_489_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_74_io_to_pes_6_out_valid = PE_490_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_74_io_to_pes_6_out_bits = PE_490_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_74_io_to_pes_7_out_valid = PE_491_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_74_io_to_pes_7_out_bits = PE_491_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_74_io_to_pes_8_out_valid = PE_492_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_74_io_to_pes_8_out_bits = PE_492_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_74_io_to_pes_9_out_valid = PE_493_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_74_io_to_pes_9_out_bits = PE_493_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_74_io_to_pes_10_out_valid = PE_494_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_74_io_to_pes_10_out_bits = PE_494_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_74_io_to_pes_11_out_valid = PE_495_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_74_io_to_pes_11_out_bits = PE_495_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_74_io_to_pes_12_out_valid = PE_496_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_74_io_to_pes_12_out_bits = PE_496_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_74_io_to_pes_13_out_valid = PE_497_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_74_io_to_pes_13_out_bits = PE_497_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_74_io_to_pes_14_out_valid = PE_498_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_74_io_to_pes_14_out_bits = PE_498_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_74_io_to_pes_15_out_valid = PE_499_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_74_io_to_pes_15_out_bits = PE_499_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_74_io_to_pes_16_out_valid = PE_500_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_74_io_to_pes_16_out_bits = PE_500_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_74_io_to_pes_17_out_valid = PE_501_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_74_io_to_pes_17_out_bits = PE_501_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_74_io_to_pes_18_out_valid = PE_502_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_74_io_to_pes_18_out_bits = PE_502_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_74_io_to_pes_19_out_valid = PE_503_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_74_io_to_pes_19_out_bits = PE_503_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_74_io_to_pes_20_out_valid = PE_504_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_74_io_to_pes_20_out_bits = PE_504_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_74_io_to_pes_21_out_valid = PE_505_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_74_io_to_pes_21_out_bits = PE_505_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_74_io_sig_stat2trans = MultiDimTime_io_index_1 == 16'h0; // @[pe.scala 278:43]
  assign PENetwork_75_clock = clock;
  assign PENetwork_75_reset = reset;
  assign PENetwork_75_io_to_pes_0_out_valid = PE_506_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_75_io_to_pes_0_out_bits = PE_506_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_75_io_to_pes_1_out_valid = PE_507_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_75_io_to_pes_1_out_bits = PE_507_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_75_io_to_pes_2_out_valid = PE_508_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_75_io_to_pes_2_out_bits = PE_508_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_75_io_to_pes_3_out_valid = PE_509_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_75_io_to_pes_3_out_bits = PE_509_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_75_io_to_pes_4_out_valid = PE_510_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_75_io_to_pes_4_out_bits = PE_510_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_75_io_to_pes_5_out_valid = PE_511_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_75_io_to_pes_5_out_bits = PE_511_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_75_io_to_pes_6_out_valid = PE_512_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_75_io_to_pes_6_out_bits = PE_512_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_75_io_to_pes_7_out_valid = PE_513_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_75_io_to_pes_7_out_bits = PE_513_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_75_io_to_pes_8_out_valid = PE_514_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_75_io_to_pes_8_out_bits = PE_514_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_75_io_to_pes_9_out_valid = PE_515_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_75_io_to_pes_9_out_bits = PE_515_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_75_io_to_pes_10_out_valid = PE_516_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_75_io_to_pes_10_out_bits = PE_516_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_75_io_to_pes_11_out_valid = PE_517_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_75_io_to_pes_11_out_bits = PE_517_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_75_io_to_pes_12_out_valid = PE_518_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_75_io_to_pes_12_out_bits = PE_518_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_75_io_to_pes_13_out_valid = PE_519_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_75_io_to_pes_13_out_bits = PE_519_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_75_io_to_pes_14_out_valid = PE_520_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_75_io_to_pes_14_out_bits = PE_520_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_75_io_to_pes_15_out_valid = PE_521_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_75_io_to_pes_15_out_bits = PE_521_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_75_io_to_pes_16_out_valid = PE_522_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_75_io_to_pes_16_out_bits = PE_522_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_75_io_to_pes_17_out_valid = PE_523_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_75_io_to_pes_17_out_bits = PE_523_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_75_io_to_pes_18_out_valid = PE_524_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_75_io_to_pes_18_out_bits = PE_524_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_75_io_to_pes_19_out_valid = PE_525_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_75_io_to_pes_19_out_bits = PE_525_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_75_io_to_pes_20_out_valid = PE_526_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_75_io_to_pes_20_out_bits = PE_526_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_75_io_to_pes_21_out_valid = PE_527_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_75_io_to_pes_21_out_bits = PE_527_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_75_io_sig_stat2trans = MultiDimTime_io_index_1 == 16'h0; // @[pe.scala 278:43]
  assign PENetwork_76_clock = clock;
  assign PENetwork_76_reset = reset;
  assign PENetwork_76_io_to_pes_0_out_valid = PE_528_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_76_io_to_pes_0_out_bits = PE_528_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_76_io_to_pes_1_out_valid = PE_529_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_76_io_to_pes_1_out_bits = PE_529_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_76_io_to_pes_2_out_valid = PE_530_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_76_io_to_pes_2_out_bits = PE_530_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_76_io_to_pes_3_out_valid = PE_531_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_76_io_to_pes_3_out_bits = PE_531_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_76_io_to_pes_4_out_valid = PE_532_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_76_io_to_pes_4_out_bits = PE_532_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_76_io_to_pes_5_out_valid = PE_533_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_76_io_to_pes_5_out_bits = PE_533_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_76_io_to_pes_6_out_valid = PE_534_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_76_io_to_pes_6_out_bits = PE_534_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_76_io_to_pes_7_out_valid = PE_535_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_76_io_to_pes_7_out_bits = PE_535_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_76_io_to_pes_8_out_valid = PE_536_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_76_io_to_pes_8_out_bits = PE_536_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_76_io_to_pes_9_out_valid = PE_537_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_76_io_to_pes_9_out_bits = PE_537_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_76_io_to_pes_10_out_valid = PE_538_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_76_io_to_pes_10_out_bits = PE_538_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_76_io_to_pes_11_out_valid = PE_539_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_76_io_to_pes_11_out_bits = PE_539_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_76_io_to_pes_12_out_valid = PE_540_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_76_io_to_pes_12_out_bits = PE_540_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_76_io_to_pes_13_out_valid = PE_541_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_76_io_to_pes_13_out_bits = PE_541_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_76_io_to_pes_14_out_valid = PE_542_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_76_io_to_pes_14_out_bits = PE_542_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_76_io_to_pes_15_out_valid = PE_543_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_76_io_to_pes_15_out_bits = PE_543_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_76_io_to_pes_16_out_valid = PE_544_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_76_io_to_pes_16_out_bits = PE_544_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_76_io_to_pes_17_out_valid = PE_545_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_76_io_to_pes_17_out_bits = PE_545_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_76_io_to_pes_18_out_valid = PE_546_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_76_io_to_pes_18_out_bits = PE_546_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_76_io_to_pes_19_out_valid = PE_547_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_76_io_to_pes_19_out_bits = PE_547_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_76_io_to_pes_20_out_valid = PE_548_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_76_io_to_pes_20_out_bits = PE_548_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_76_io_to_pes_21_out_valid = PE_549_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_76_io_to_pes_21_out_bits = PE_549_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_76_io_sig_stat2trans = MultiDimTime_io_index_1 == 16'h0; // @[pe.scala 278:43]
  assign PENetwork_77_clock = clock;
  assign PENetwork_77_reset = reset;
  assign PENetwork_77_io_to_pes_0_out_valid = PE_550_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_77_io_to_pes_0_out_bits = PE_550_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_77_io_to_pes_1_out_valid = PE_551_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_77_io_to_pes_1_out_bits = PE_551_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_77_io_to_pes_2_out_valid = PE_552_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_77_io_to_pes_2_out_bits = PE_552_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_77_io_to_pes_3_out_valid = PE_553_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_77_io_to_pes_3_out_bits = PE_553_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_77_io_to_pes_4_out_valid = PE_554_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_77_io_to_pes_4_out_bits = PE_554_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_77_io_to_pes_5_out_valid = PE_555_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_77_io_to_pes_5_out_bits = PE_555_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_77_io_to_pes_6_out_valid = PE_556_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_77_io_to_pes_6_out_bits = PE_556_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_77_io_to_pes_7_out_valid = PE_557_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_77_io_to_pes_7_out_bits = PE_557_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_77_io_to_pes_8_out_valid = PE_558_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_77_io_to_pes_8_out_bits = PE_558_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_77_io_to_pes_9_out_valid = PE_559_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_77_io_to_pes_9_out_bits = PE_559_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_77_io_to_pes_10_out_valid = PE_560_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_77_io_to_pes_10_out_bits = PE_560_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_77_io_to_pes_11_out_valid = PE_561_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_77_io_to_pes_11_out_bits = PE_561_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_77_io_to_pes_12_out_valid = PE_562_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_77_io_to_pes_12_out_bits = PE_562_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_77_io_to_pes_13_out_valid = PE_563_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_77_io_to_pes_13_out_bits = PE_563_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_77_io_to_pes_14_out_valid = PE_564_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_77_io_to_pes_14_out_bits = PE_564_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_77_io_to_pes_15_out_valid = PE_565_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_77_io_to_pes_15_out_bits = PE_565_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_77_io_to_pes_16_out_valid = PE_566_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_77_io_to_pes_16_out_bits = PE_566_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_77_io_to_pes_17_out_valid = PE_567_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_77_io_to_pes_17_out_bits = PE_567_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_77_io_to_pes_18_out_valid = PE_568_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_77_io_to_pes_18_out_bits = PE_568_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_77_io_to_pes_19_out_valid = PE_569_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_77_io_to_pes_19_out_bits = PE_569_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_77_io_to_pes_20_out_valid = PE_570_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_77_io_to_pes_20_out_bits = PE_570_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_77_io_to_pes_21_out_valid = PE_571_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_77_io_to_pes_21_out_bits = PE_571_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_77_io_sig_stat2trans = MultiDimTime_io_index_1 == 16'h0; // @[pe.scala 278:43]
  assign PENetwork_78_clock = clock;
  assign PENetwork_78_reset = reset;
  assign PENetwork_78_io_to_pes_0_out_valid = PE_572_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_78_io_to_pes_0_out_bits = PE_572_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_78_io_to_pes_1_out_valid = PE_573_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_78_io_to_pes_1_out_bits = PE_573_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_78_io_to_pes_2_out_valid = PE_574_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_78_io_to_pes_2_out_bits = PE_574_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_78_io_to_pes_3_out_valid = PE_575_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_78_io_to_pes_3_out_bits = PE_575_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_78_io_to_pes_4_out_valid = PE_576_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_78_io_to_pes_4_out_bits = PE_576_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_78_io_to_pes_5_out_valid = PE_577_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_78_io_to_pes_5_out_bits = PE_577_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_78_io_to_pes_6_out_valid = PE_578_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_78_io_to_pes_6_out_bits = PE_578_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_78_io_to_pes_7_out_valid = PE_579_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_78_io_to_pes_7_out_bits = PE_579_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_78_io_to_pes_8_out_valid = PE_580_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_78_io_to_pes_8_out_bits = PE_580_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_78_io_to_pes_9_out_valid = PE_581_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_78_io_to_pes_9_out_bits = PE_581_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_78_io_to_pes_10_out_valid = PE_582_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_78_io_to_pes_10_out_bits = PE_582_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_78_io_to_pes_11_out_valid = PE_583_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_78_io_to_pes_11_out_bits = PE_583_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_78_io_to_pes_12_out_valid = PE_584_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_78_io_to_pes_12_out_bits = PE_584_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_78_io_to_pes_13_out_valid = PE_585_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_78_io_to_pes_13_out_bits = PE_585_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_78_io_to_pes_14_out_valid = PE_586_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_78_io_to_pes_14_out_bits = PE_586_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_78_io_to_pes_15_out_valid = PE_587_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_78_io_to_pes_15_out_bits = PE_587_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_78_io_to_pes_16_out_valid = PE_588_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_78_io_to_pes_16_out_bits = PE_588_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_78_io_to_pes_17_out_valid = PE_589_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_78_io_to_pes_17_out_bits = PE_589_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_78_io_to_pes_18_out_valid = PE_590_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_78_io_to_pes_18_out_bits = PE_590_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_78_io_to_pes_19_out_valid = PE_591_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_78_io_to_pes_19_out_bits = PE_591_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_78_io_to_pes_20_out_valid = PE_592_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_78_io_to_pes_20_out_bits = PE_592_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_78_io_to_pes_21_out_valid = PE_593_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_78_io_to_pes_21_out_bits = PE_593_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_78_io_sig_stat2trans = MultiDimTime_io_index_1 == 16'h0; // @[pe.scala 278:43]
  assign PENetwork_79_clock = clock;
  assign PENetwork_79_reset = reset;
  assign PENetwork_79_io_to_pes_0_out_valid = PE_594_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_79_io_to_pes_0_out_bits = PE_594_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_79_io_to_pes_1_out_valid = PE_595_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_79_io_to_pes_1_out_bits = PE_595_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_79_io_to_pes_2_out_valid = PE_596_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_79_io_to_pes_2_out_bits = PE_596_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_79_io_to_pes_3_out_valid = PE_597_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_79_io_to_pes_3_out_bits = PE_597_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_79_io_to_pes_4_out_valid = PE_598_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_79_io_to_pes_4_out_bits = PE_598_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_79_io_to_pes_5_out_valid = PE_599_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_79_io_to_pes_5_out_bits = PE_599_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_79_io_to_pes_6_out_valid = PE_600_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_79_io_to_pes_6_out_bits = PE_600_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_79_io_to_pes_7_out_valid = PE_601_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_79_io_to_pes_7_out_bits = PE_601_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_79_io_to_pes_8_out_valid = PE_602_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_79_io_to_pes_8_out_bits = PE_602_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_79_io_to_pes_9_out_valid = PE_603_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_79_io_to_pes_9_out_bits = PE_603_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_79_io_to_pes_10_out_valid = PE_604_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_79_io_to_pes_10_out_bits = PE_604_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_79_io_to_pes_11_out_valid = PE_605_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_79_io_to_pes_11_out_bits = PE_605_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_79_io_to_pes_12_out_valid = PE_606_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_79_io_to_pes_12_out_bits = PE_606_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_79_io_to_pes_13_out_valid = PE_607_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_79_io_to_pes_13_out_bits = PE_607_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_79_io_to_pes_14_out_valid = PE_608_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_79_io_to_pes_14_out_bits = PE_608_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_79_io_to_pes_15_out_valid = PE_609_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_79_io_to_pes_15_out_bits = PE_609_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_79_io_to_pes_16_out_valid = PE_610_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_79_io_to_pes_16_out_bits = PE_610_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_79_io_to_pes_17_out_valid = PE_611_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_79_io_to_pes_17_out_bits = PE_611_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_79_io_to_pes_18_out_valid = PE_612_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_79_io_to_pes_18_out_bits = PE_612_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_79_io_to_pes_19_out_valid = PE_613_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_79_io_to_pes_19_out_bits = PE_613_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_79_io_to_pes_20_out_valid = PE_614_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_79_io_to_pes_20_out_bits = PE_614_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_79_io_to_pes_21_out_valid = PE_615_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_79_io_to_pes_21_out_bits = PE_615_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_79_io_sig_stat2trans = MultiDimTime_io_index_1 == 16'h0; // @[pe.scala 278:43]
  assign PENetwork_80_clock = clock;
  assign PENetwork_80_reset = reset;
  assign PENetwork_80_io_to_pes_0_out_valid = PE_616_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_80_io_to_pes_0_out_bits = PE_616_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_80_io_to_pes_1_out_valid = PE_617_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_80_io_to_pes_1_out_bits = PE_617_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_80_io_to_pes_2_out_valid = PE_618_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_80_io_to_pes_2_out_bits = PE_618_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_80_io_to_pes_3_out_valid = PE_619_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_80_io_to_pes_3_out_bits = PE_619_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_80_io_to_pes_4_out_valid = PE_620_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_80_io_to_pes_4_out_bits = PE_620_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_80_io_to_pes_5_out_valid = PE_621_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_80_io_to_pes_5_out_bits = PE_621_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_80_io_to_pes_6_out_valid = PE_622_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_80_io_to_pes_6_out_bits = PE_622_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_80_io_to_pes_7_out_valid = PE_623_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_80_io_to_pes_7_out_bits = PE_623_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_80_io_to_pes_8_out_valid = PE_624_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_80_io_to_pes_8_out_bits = PE_624_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_80_io_to_pes_9_out_valid = PE_625_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_80_io_to_pes_9_out_bits = PE_625_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_80_io_to_pes_10_out_valid = PE_626_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_80_io_to_pes_10_out_bits = PE_626_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_80_io_to_pes_11_out_valid = PE_627_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_80_io_to_pes_11_out_bits = PE_627_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_80_io_to_pes_12_out_valid = PE_628_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_80_io_to_pes_12_out_bits = PE_628_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_80_io_to_pes_13_out_valid = PE_629_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_80_io_to_pes_13_out_bits = PE_629_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_80_io_to_pes_14_out_valid = PE_630_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_80_io_to_pes_14_out_bits = PE_630_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_80_io_to_pes_15_out_valid = PE_631_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_80_io_to_pes_15_out_bits = PE_631_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_80_io_to_pes_16_out_valid = PE_632_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_80_io_to_pes_16_out_bits = PE_632_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_80_io_to_pes_17_out_valid = PE_633_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_80_io_to_pes_17_out_bits = PE_633_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_80_io_to_pes_18_out_valid = PE_634_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_80_io_to_pes_18_out_bits = PE_634_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_80_io_to_pes_19_out_valid = PE_635_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_80_io_to_pes_19_out_bits = PE_635_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_80_io_to_pes_20_out_valid = PE_636_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_80_io_to_pes_20_out_bits = PE_636_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_80_io_to_pes_21_out_valid = PE_637_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_80_io_to_pes_21_out_bits = PE_637_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_80_io_sig_stat2trans = MultiDimTime_io_index_1 == 16'h0; // @[pe.scala 278:43]
  assign PENetwork_81_clock = clock;
  assign PENetwork_81_reset = reset;
  assign PENetwork_81_io_to_pes_0_out_valid = PE_638_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_81_io_to_pes_0_out_bits = PE_638_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_81_io_to_pes_1_out_valid = PE_639_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_81_io_to_pes_1_out_bits = PE_639_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_81_io_to_pes_2_out_valid = PE_640_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_81_io_to_pes_2_out_bits = PE_640_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_81_io_to_pes_3_out_valid = PE_641_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_81_io_to_pes_3_out_bits = PE_641_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_81_io_to_pes_4_out_valid = PE_642_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_81_io_to_pes_4_out_bits = PE_642_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_81_io_to_pes_5_out_valid = PE_643_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_81_io_to_pes_5_out_bits = PE_643_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_81_io_to_pes_6_out_valid = PE_644_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_81_io_to_pes_6_out_bits = PE_644_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_81_io_to_pes_7_out_valid = PE_645_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_81_io_to_pes_7_out_bits = PE_645_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_81_io_to_pes_8_out_valid = PE_646_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_81_io_to_pes_8_out_bits = PE_646_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_81_io_to_pes_9_out_valid = PE_647_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_81_io_to_pes_9_out_bits = PE_647_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_81_io_to_pes_10_out_valid = PE_648_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_81_io_to_pes_10_out_bits = PE_648_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_81_io_to_pes_11_out_valid = PE_649_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_81_io_to_pes_11_out_bits = PE_649_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_81_io_to_pes_12_out_valid = PE_650_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_81_io_to_pes_12_out_bits = PE_650_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_81_io_to_pes_13_out_valid = PE_651_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_81_io_to_pes_13_out_bits = PE_651_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_81_io_to_pes_14_out_valid = PE_652_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_81_io_to_pes_14_out_bits = PE_652_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_81_io_to_pes_15_out_valid = PE_653_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_81_io_to_pes_15_out_bits = PE_653_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_81_io_to_pes_16_out_valid = PE_654_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_81_io_to_pes_16_out_bits = PE_654_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_81_io_to_pes_17_out_valid = PE_655_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_81_io_to_pes_17_out_bits = PE_655_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_81_io_to_pes_18_out_valid = PE_656_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_81_io_to_pes_18_out_bits = PE_656_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_81_io_to_pes_19_out_valid = PE_657_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_81_io_to_pes_19_out_bits = PE_657_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_81_io_to_pes_20_out_valid = PE_658_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_81_io_to_pes_20_out_bits = PE_658_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_81_io_to_pes_21_out_valid = PE_659_io_data_2_out_valid; // @[pe.scala 263:36]
  assign PENetwork_81_io_to_pes_21_out_bits = PE_659_io_data_2_out_bits; // @[pe.scala 263:36]
  assign PENetwork_81_io_sig_stat2trans = MultiDimTime_io_index_1 == 16'h0; // @[pe.scala 278:43]
  assign MemController_clock = clock;
  assign MemController_reset = reset;
  assign MemController_io_rd_valid = io_exec_valid; // @[pe.scala 310:28]
  assign MemController_io_wr_valid = io_data_0_in_0_valid; // @[pe.scala 311:28]
  assign MemController_io_wr_data_valid = io_data_0_in_0_bits_valid; // @[pe.scala 313:27]
  assign MemController_io_wr_data_bits = io_data_0_in_0_bits_bits; // @[pe.scala 313:27]
  assign MemController_1_clock = clock;
  assign MemController_1_reset = reset;
  assign MemController_1_io_rd_valid = io_exec_valid; // @[pe.scala 310:28]
  assign MemController_1_io_wr_valid = io_data_0_in_1_valid; // @[pe.scala 311:28]
  assign MemController_1_io_wr_data_valid = io_data_0_in_1_bits_valid; // @[pe.scala 313:27]
  assign MemController_1_io_wr_data_bits = io_data_0_in_1_bits_bits; // @[pe.scala 313:27]
  assign MemController_2_clock = clock;
  assign MemController_2_reset = reset;
  assign MemController_2_io_rd_valid = io_exec_valid; // @[pe.scala 310:28]
  assign MemController_2_io_wr_valid = io_data_0_in_2_valid; // @[pe.scala 311:28]
  assign MemController_2_io_wr_data_valid = io_data_0_in_2_bits_valid; // @[pe.scala 313:27]
  assign MemController_2_io_wr_data_bits = io_data_0_in_2_bits_bits; // @[pe.scala 313:27]
  assign MemController_3_clock = clock;
  assign MemController_3_reset = reset;
  assign MemController_3_io_rd_valid = io_exec_valid; // @[pe.scala 310:28]
  assign MemController_3_io_wr_valid = io_data_0_in_3_valid; // @[pe.scala 311:28]
  assign MemController_3_io_wr_data_valid = io_data_0_in_3_bits_valid; // @[pe.scala 313:27]
  assign MemController_3_io_wr_data_bits = io_data_0_in_3_bits_bits; // @[pe.scala 313:27]
  assign MemController_4_clock = clock;
  assign MemController_4_reset = reset;
  assign MemController_4_io_rd_valid = io_exec_valid; // @[pe.scala 310:28]
  assign MemController_4_io_wr_valid = io_data_0_in_4_valid; // @[pe.scala 311:28]
  assign MemController_4_io_wr_data_valid = io_data_0_in_4_bits_valid; // @[pe.scala 313:27]
  assign MemController_4_io_wr_data_bits = io_data_0_in_4_bits_bits; // @[pe.scala 313:27]
  assign MemController_5_clock = clock;
  assign MemController_5_reset = reset;
  assign MemController_5_io_rd_valid = io_exec_valid; // @[pe.scala 310:28]
  assign MemController_5_io_wr_valid = io_data_0_in_5_valid; // @[pe.scala 311:28]
  assign MemController_5_io_wr_data_valid = io_data_0_in_5_bits_valid; // @[pe.scala 313:27]
  assign MemController_5_io_wr_data_bits = io_data_0_in_5_bits_bits; // @[pe.scala 313:27]
  assign MemController_6_clock = clock;
  assign MemController_6_reset = reset;
  assign MemController_6_io_rd_valid = io_exec_valid; // @[pe.scala 310:28]
  assign MemController_6_io_wr_valid = io_data_0_in_6_valid; // @[pe.scala 311:28]
  assign MemController_6_io_wr_data_valid = io_data_0_in_6_bits_valid; // @[pe.scala 313:27]
  assign MemController_6_io_wr_data_bits = io_data_0_in_6_bits_bits; // @[pe.scala 313:27]
  assign MemController_7_clock = clock;
  assign MemController_7_reset = reset;
  assign MemController_7_io_rd_valid = io_exec_valid; // @[pe.scala 310:28]
  assign MemController_7_io_wr_valid = io_data_0_in_7_valid; // @[pe.scala 311:28]
  assign MemController_7_io_wr_data_valid = io_data_0_in_7_bits_valid; // @[pe.scala 313:27]
  assign MemController_7_io_wr_data_bits = io_data_0_in_7_bits_bits; // @[pe.scala 313:27]
  assign MemController_8_clock = clock;
  assign MemController_8_reset = reset;
  assign MemController_8_io_rd_valid = io_exec_valid; // @[pe.scala 310:28]
  assign MemController_8_io_wr_valid = io_data_0_in_8_valid; // @[pe.scala 311:28]
  assign MemController_8_io_wr_data_valid = io_data_0_in_8_bits_valid; // @[pe.scala 313:27]
  assign MemController_8_io_wr_data_bits = io_data_0_in_8_bits_bits; // @[pe.scala 313:27]
  assign MemController_9_clock = clock;
  assign MemController_9_reset = reset;
  assign MemController_9_io_rd_valid = io_exec_valid; // @[pe.scala 310:28]
  assign MemController_9_io_wr_valid = io_data_0_in_9_valid; // @[pe.scala 311:28]
  assign MemController_9_io_wr_data_valid = io_data_0_in_9_bits_valid; // @[pe.scala 313:27]
  assign MemController_9_io_wr_data_bits = io_data_0_in_9_bits_bits; // @[pe.scala 313:27]
  assign MemController_10_clock = clock;
  assign MemController_10_reset = reset;
  assign MemController_10_io_rd_valid = io_exec_valid; // @[pe.scala 310:28]
  assign MemController_10_io_wr_valid = io_data_0_in_10_valid; // @[pe.scala 311:28]
  assign MemController_10_io_wr_data_valid = io_data_0_in_10_bits_valid; // @[pe.scala 313:27]
  assign MemController_10_io_wr_data_bits = io_data_0_in_10_bits_bits; // @[pe.scala 313:27]
  assign MemController_11_clock = clock;
  assign MemController_11_reset = reset;
  assign MemController_11_io_rd_valid = io_exec_valid; // @[pe.scala 310:28]
  assign MemController_11_io_wr_valid = io_data_0_in_11_valid; // @[pe.scala 311:28]
  assign MemController_11_io_wr_data_valid = io_data_0_in_11_bits_valid; // @[pe.scala 313:27]
  assign MemController_11_io_wr_data_bits = io_data_0_in_11_bits_bits; // @[pe.scala 313:27]
  assign MemController_12_clock = clock;
  assign MemController_12_reset = reset;
  assign MemController_12_io_rd_valid = io_exec_valid; // @[pe.scala 310:28]
  assign MemController_12_io_wr_valid = io_data_0_in_12_valid; // @[pe.scala 311:28]
  assign MemController_12_io_wr_data_valid = io_data_0_in_12_bits_valid; // @[pe.scala 313:27]
  assign MemController_12_io_wr_data_bits = io_data_0_in_12_bits_bits; // @[pe.scala 313:27]
  assign MemController_13_clock = clock;
  assign MemController_13_reset = reset;
  assign MemController_13_io_rd_valid = io_exec_valid; // @[pe.scala 310:28]
  assign MemController_13_io_wr_valid = io_data_0_in_13_valid; // @[pe.scala 311:28]
  assign MemController_13_io_wr_data_valid = io_data_0_in_13_bits_valid; // @[pe.scala 313:27]
  assign MemController_13_io_wr_data_bits = io_data_0_in_13_bits_bits; // @[pe.scala 313:27]
  assign MemController_14_clock = clock;
  assign MemController_14_reset = reset;
  assign MemController_14_io_rd_valid = io_exec_valid; // @[pe.scala 310:28]
  assign MemController_14_io_wr_valid = io_data_0_in_14_valid; // @[pe.scala 311:28]
  assign MemController_14_io_wr_data_valid = io_data_0_in_14_bits_valid; // @[pe.scala 313:27]
  assign MemController_14_io_wr_data_bits = io_data_0_in_14_bits_bits; // @[pe.scala 313:27]
  assign MemController_15_clock = clock;
  assign MemController_15_reset = reset;
  assign MemController_15_io_rd_valid = io_exec_valid; // @[pe.scala 310:28]
  assign MemController_15_io_wr_valid = io_data_0_in_15_valid; // @[pe.scala 311:28]
  assign MemController_15_io_wr_data_valid = io_data_0_in_15_bits_valid; // @[pe.scala 313:27]
  assign MemController_15_io_wr_data_bits = io_data_0_in_15_bits_bits; // @[pe.scala 313:27]
  assign MemController_16_clock = clock;
  assign MemController_16_reset = reset;
  assign MemController_16_io_rd_valid = io_exec_valid; // @[pe.scala 310:28]
  assign MemController_16_io_wr_valid = io_data_0_in_16_valid; // @[pe.scala 311:28]
  assign MemController_16_io_wr_data_valid = io_data_0_in_16_bits_valid; // @[pe.scala 313:27]
  assign MemController_16_io_wr_data_bits = io_data_0_in_16_bits_bits; // @[pe.scala 313:27]
  assign MemController_17_clock = clock;
  assign MemController_17_reset = reset;
  assign MemController_17_io_rd_valid = io_exec_valid; // @[pe.scala 310:28]
  assign MemController_17_io_wr_valid = io_data_0_in_17_valid; // @[pe.scala 311:28]
  assign MemController_17_io_wr_data_valid = io_data_0_in_17_bits_valid; // @[pe.scala 313:27]
  assign MemController_17_io_wr_data_bits = io_data_0_in_17_bits_bits; // @[pe.scala 313:27]
  assign MemController_18_clock = clock;
  assign MemController_18_reset = reset;
  assign MemController_18_io_rd_valid = io_exec_valid; // @[pe.scala 310:28]
  assign MemController_18_io_wr_valid = io_data_0_in_18_valid; // @[pe.scala 311:28]
  assign MemController_18_io_wr_data_valid = io_data_0_in_18_bits_valid; // @[pe.scala 313:27]
  assign MemController_18_io_wr_data_bits = io_data_0_in_18_bits_bits; // @[pe.scala 313:27]
  assign MemController_19_clock = clock;
  assign MemController_19_reset = reset;
  assign MemController_19_io_rd_valid = io_exec_valid; // @[pe.scala 310:28]
  assign MemController_19_io_wr_valid = io_data_0_in_19_valid; // @[pe.scala 311:28]
  assign MemController_19_io_wr_data_valid = io_data_0_in_19_bits_valid; // @[pe.scala 313:27]
  assign MemController_19_io_wr_data_bits = io_data_0_in_19_bits_bits; // @[pe.scala 313:27]
  assign MemController_20_clock = clock;
  assign MemController_20_reset = reset;
  assign MemController_20_io_rd_valid = io_exec_valid; // @[pe.scala 310:28]
  assign MemController_20_io_wr_valid = io_data_0_in_20_valid; // @[pe.scala 311:28]
  assign MemController_20_io_wr_data_valid = io_data_0_in_20_bits_valid; // @[pe.scala 313:27]
  assign MemController_20_io_wr_data_bits = io_data_0_in_20_bits_bits; // @[pe.scala 313:27]
  assign MemController_21_clock = clock;
  assign MemController_21_reset = reset;
  assign MemController_21_io_rd_valid = io_exec_valid; // @[pe.scala 310:28]
  assign MemController_21_io_wr_valid = io_data_0_in_21_valid; // @[pe.scala 311:28]
  assign MemController_21_io_wr_data_valid = io_data_0_in_21_bits_valid; // @[pe.scala 313:27]
  assign MemController_21_io_wr_data_bits = io_data_0_in_21_bits_bits; // @[pe.scala 313:27]
  assign MemController_22_clock = clock;
  assign MemController_22_reset = reset;
  assign MemController_22_io_rd_valid = io_exec_valid; // @[pe.scala 310:28]
  assign MemController_22_io_wr_valid = io_data_1_in_0_valid; // @[pe.scala 311:28]
  assign MemController_22_io_wr_data_valid = io_data_1_in_0_bits_valid; // @[pe.scala 313:27]
  assign MemController_22_io_wr_data_bits = io_data_1_in_0_bits_bits; // @[pe.scala 313:27]
  assign MemController_23_clock = clock;
  assign MemController_23_reset = reset;
  assign MemController_23_io_rd_valid = io_exec_valid; // @[pe.scala 310:28]
  assign MemController_23_io_wr_valid = io_data_1_in_1_valid; // @[pe.scala 311:28]
  assign MemController_23_io_wr_data_valid = io_data_1_in_1_bits_valid; // @[pe.scala 313:27]
  assign MemController_23_io_wr_data_bits = io_data_1_in_1_bits_bits; // @[pe.scala 313:27]
  assign MemController_24_clock = clock;
  assign MemController_24_reset = reset;
  assign MemController_24_io_rd_valid = io_exec_valid; // @[pe.scala 310:28]
  assign MemController_24_io_wr_valid = io_data_1_in_2_valid; // @[pe.scala 311:28]
  assign MemController_24_io_wr_data_valid = io_data_1_in_2_bits_valid; // @[pe.scala 313:27]
  assign MemController_24_io_wr_data_bits = io_data_1_in_2_bits_bits; // @[pe.scala 313:27]
  assign MemController_25_clock = clock;
  assign MemController_25_reset = reset;
  assign MemController_25_io_rd_valid = io_exec_valid; // @[pe.scala 310:28]
  assign MemController_25_io_wr_valid = io_data_1_in_3_valid; // @[pe.scala 311:28]
  assign MemController_25_io_wr_data_valid = io_data_1_in_3_bits_valid; // @[pe.scala 313:27]
  assign MemController_25_io_wr_data_bits = io_data_1_in_3_bits_bits; // @[pe.scala 313:27]
  assign MemController_26_clock = clock;
  assign MemController_26_reset = reset;
  assign MemController_26_io_rd_valid = io_exec_valid; // @[pe.scala 310:28]
  assign MemController_26_io_wr_valid = io_data_1_in_4_valid; // @[pe.scala 311:28]
  assign MemController_26_io_wr_data_valid = io_data_1_in_4_bits_valid; // @[pe.scala 313:27]
  assign MemController_26_io_wr_data_bits = io_data_1_in_4_bits_bits; // @[pe.scala 313:27]
  assign MemController_27_clock = clock;
  assign MemController_27_reset = reset;
  assign MemController_27_io_rd_valid = io_exec_valid; // @[pe.scala 310:28]
  assign MemController_27_io_wr_valid = io_data_1_in_5_valid; // @[pe.scala 311:28]
  assign MemController_27_io_wr_data_valid = io_data_1_in_5_bits_valid; // @[pe.scala 313:27]
  assign MemController_27_io_wr_data_bits = io_data_1_in_5_bits_bits; // @[pe.scala 313:27]
  assign MemController_28_clock = clock;
  assign MemController_28_reset = reset;
  assign MemController_28_io_rd_valid = io_exec_valid; // @[pe.scala 310:28]
  assign MemController_28_io_wr_valid = io_data_1_in_6_valid; // @[pe.scala 311:28]
  assign MemController_28_io_wr_data_valid = io_data_1_in_6_bits_valid; // @[pe.scala 313:27]
  assign MemController_28_io_wr_data_bits = io_data_1_in_6_bits_bits; // @[pe.scala 313:27]
  assign MemController_29_clock = clock;
  assign MemController_29_reset = reset;
  assign MemController_29_io_rd_valid = io_exec_valid; // @[pe.scala 310:28]
  assign MemController_29_io_wr_valid = io_data_1_in_7_valid; // @[pe.scala 311:28]
  assign MemController_29_io_wr_data_valid = io_data_1_in_7_bits_valid; // @[pe.scala 313:27]
  assign MemController_29_io_wr_data_bits = io_data_1_in_7_bits_bits; // @[pe.scala 313:27]
  assign MemController_30_clock = clock;
  assign MemController_30_reset = reset;
  assign MemController_30_io_rd_valid = io_exec_valid; // @[pe.scala 310:28]
  assign MemController_30_io_wr_valid = io_data_1_in_8_valid; // @[pe.scala 311:28]
  assign MemController_30_io_wr_data_valid = io_data_1_in_8_bits_valid; // @[pe.scala 313:27]
  assign MemController_30_io_wr_data_bits = io_data_1_in_8_bits_bits; // @[pe.scala 313:27]
  assign MemController_31_clock = clock;
  assign MemController_31_reset = reset;
  assign MemController_31_io_rd_valid = io_exec_valid; // @[pe.scala 310:28]
  assign MemController_31_io_wr_valid = io_data_1_in_9_valid; // @[pe.scala 311:28]
  assign MemController_31_io_wr_data_valid = io_data_1_in_9_bits_valid; // @[pe.scala 313:27]
  assign MemController_31_io_wr_data_bits = io_data_1_in_9_bits_bits; // @[pe.scala 313:27]
  assign MemController_32_clock = clock;
  assign MemController_32_reset = reset;
  assign MemController_32_io_rd_valid = io_exec_valid; // @[pe.scala 310:28]
  assign MemController_32_io_wr_valid = io_data_1_in_10_valid; // @[pe.scala 311:28]
  assign MemController_32_io_wr_data_valid = io_data_1_in_10_bits_valid; // @[pe.scala 313:27]
  assign MemController_32_io_wr_data_bits = io_data_1_in_10_bits_bits; // @[pe.scala 313:27]
  assign MemController_33_clock = clock;
  assign MemController_33_reset = reset;
  assign MemController_33_io_rd_valid = io_exec_valid; // @[pe.scala 310:28]
  assign MemController_33_io_wr_valid = io_data_1_in_11_valid; // @[pe.scala 311:28]
  assign MemController_33_io_wr_data_valid = io_data_1_in_11_bits_valid; // @[pe.scala 313:27]
  assign MemController_33_io_wr_data_bits = io_data_1_in_11_bits_bits; // @[pe.scala 313:27]
  assign MemController_34_clock = clock;
  assign MemController_34_reset = reset;
  assign MemController_34_io_rd_valid = io_exec_valid; // @[pe.scala 310:28]
  assign MemController_34_io_wr_valid = io_data_1_in_12_valid; // @[pe.scala 311:28]
  assign MemController_34_io_wr_data_valid = io_data_1_in_12_bits_valid; // @[pe.scala 313:27]
  assign MemController_34_io_wr_data_bits = io_data_1_in_12_bits_bits; // @[pe.scala 313:27]
  assign MemController_35_clock = clock;
  assign MemController_35_reset = reset;
  assign MemController_35_io_rd_valid = io_exec_valid; // @[pe.scala 310:28]
  assign MemController_35_io_wr_valid = io_data_1_in_13_valid; // @[pe.scala 311:28]
  assign MemController_35_io_wr_data_valid = io_data_1_in_13_bits_valid; // @[pe.scala 313:27]
  assign MemController_35_io_wr_data_bits = io_data_1_in_13_bits_bits; // @[pe.scala 313:27]
  assign MemController_36_clock = clock;
  assign MemController_36_reset = reset;
  assign MemController_36_io_rd_valid = io_exec_valid; // @[pe.scala 310:28]
  assign MemController_36_io_wr_valid = io_data_1_in_14_valid; // @[pe.scala 311:28]
  assign MemController_36_io_wr_data_valid = io_data_1_in_14_bits_valid; // @[pe.scala 313:27]
  assign MemController_36_io_wr_data_bits = io_data_1_in_14_bits_bits; // @[pe.scala 313:27]
  assign MemController_37_clock = clock;
  assign MemController_37_reset = reset;
  assign MemController_37_io_rd_valid = io_exec_valid; // @[pe.scala 310:28]
  assign MemController_37_io_wr_valid = io_data_1_in_15_valid; // @[pe.scala 311:28]
  assign MemController_37_io_wr_data_valid = io_data_1_in_15_bits_valid; // @[pe.scala 313:27]
  assign MemController_37_io_wr_data_bits = io_data_1_in_15_bits_bits; // @[pe.scala 313:27]
  assign MemController_38_clock = clock;
  assign MemController_38_reset = reset;
  assign MemController_38_io_rd_valid = io_exec_valid; // @[pe.scala 310:28]
  assign MemController_38_io_wr_valid = io_data_1_in_16_valid; // @[pe.scala 311:28]
  assign MemController_38_io_wr_data_valid = io_data_1_in_16_bits_valid; // @[pe.scala 313:27]
  assign MemController_38_io_wr_data_bits = io_data_1_in_16_bits_bits; // @[pe.scala 313:27]
  assign MemController_39_clock = clock;
  assign MemController_39_reset = reset;
  assign MemController_39_io_rd_valid = io_exec_valid; // @[pe.scala 310:28]
  assign MemController_39_io_wr_valid = io_data_1_in_17_valid; // @[pe.scala 311:28]
  assign MemController_39_io_wr_data_valid = io_data_1_in_17_bits_valid; // @[pe.scala 313:27]
  assign MemController_39_io_wr_data_bits = io_data_1_in_17_bits_bits; // @[pe.scala 313:27]
  assign MemController_40_clock = clock;
  assign MemController_40_reset = reset;
  assign MemController_40_io_rd_valid = io_exec_valid; // @[pe.scala 310:28]
  assign MemController_40_io_wr_valid = io_data_1_in_18_valid; // @[pe.scala 311:28]
  assign MemController_40_io_wr_data_valid = io_data_1_in_18_bits_valid; // @[pe.scala 313:27]
  assign MemController_40_io_wr_data_bits = io_data_1_in_18_bits_bits; // @[pe.scala 313:27]
  assign MemController_41_clock = clock;
  assign MemController_41_reset = reset;
  assign MemController_41_io_rd_valid = io_exec_valid; // @[pe.scala 310:28]
  assign MemController_41_io_wr_valid = io_data_1_in_19_valid; // @[pe.scala 311:28]
  assign MemController_41_io_wr_data_valid = io_data_1_in_19_bits_valid; // @[pe.scala 313:27]
  assign MemController_41_io_wr_data_bits = io_data_1_in_19_bits_bits; // @[pe.scala 313:27]
  assign MemController_42_clock = clock;
  assign MemController_42_reset = reset;
  assign MemController_42_io_rd_valid = io_exec_valid; // @[pe.scala 310:28]
  assign MemController_42_io_wr_valid = io_data_1_in_20_valid; // @[pe.scala 311:28]
  assign MemController_42_io_wr_data_valid = io_data_1_in_20_bits_valid; // @[pe.scala 313:27]
  assign MemController_42_io_wr_data_bits = io_data_1_in_20_bits_bits; // @[pe.scala 313:27]
  assign MemController_43_clock = clock;
  assign MemController_43_reset = reset;
  assign MemController_43_io_rd_valid = io_exec_valid; // @[pe.scala 310:28]
  assign MemController_43_io_wr_valid = io_data_1_in_21_valid; // @[pe.scala 311:28]
  assign MemController_43_io_wr_data_valid = io_data_1_in_21_bits_valid; // @[pe.scala 313:27]
  assign MemController_43_io_wr_data_bits = io_data_1_in_21_bits_bits; // @[pe.scala 313:27]
  assign MemController_44_clock = clock;
  assign MemController_44_reset = reset;
  assign MemController_44_io_rd_valid = io_exec_valid; // @[pe.scala 310:28]
  assign MemController_44_io_wr_valid = io_data_1_in_22_valid; // @[pe.scala 311:28]
  assign MemController_44_io_wr_data_valid = io_data_1_in_22_bits_valid; // @[pe.scala 313:27]
  assign MemController_44_io_wr_data_bits = io_data_1_in_22_bits_bits; // @[pe.scala 313:27]
  assign MemController_45_clock = clock;
  assign MemController_45_reset = reset;
  assign MemController_45_io_rd_valid = io_exec_valid; // @[pe.scala 310:28]
  assign MemController_45_io_wr_valid = io_data_1_in_23_valid; // @[pe.scala 311:28]
  assign MemController_45_io_wr_data_valid = io_data_1_in_23_bits_valid; // @[pe.scala 313:27]
  assign MemController_45_io_wr_data_bits = io_data_1_in_23_bits_bits; // @[pe.scala 313:27]
  assign MemController_46_clock = clock;
  assign MemController_46_reset = reset;
  assign MemController_46_io_rd_valid = io_exec_valid; // @[pe.scala 310:28]
  assign MemController_46_io_wr_valid = io_data_1_in_24_valid; // @[pe.scala 311:28]
  assign MemController_46_io_wr_data_valid = io_data_1_in_24_bits_valid; // @[pe.scala 313:27]
  assign MemController_46_io_wr_data_bits = io_data_1_in_24_bits_bits; // @[pe.scala 313:27]
  assign MemController_47_clock = clock;
  assign MemController_47_reset = reset;
  assign MemController_47_io_rd_valid = io_exec_valid; // @[pe.scala 310:28]
  assign MemController_47_io_wr_valid = io_data_1_in_25_valid; // @[pe.scala 311:28]
  assign MemController_47_io_wr_data_valid = io_data_1_in_25_bits_valid; // @[pe.scala 313:27]
  assign MemController_47_io_wr_data_bits = io_data_1_in_25_bits_bits; // @[pe.scala 313:27]
  assign MemController_48_clock = clock;
  assign MemController_48_reset = reset;
  assign MemController_48_io_rd_valid = io_exec_valid; // @[pe.scala 310:28]
  assign MemController_48_io_wr_valid = io_data_1_in_26_valid; // @[pe.scala 311:28]
  assign MemController_48_io_wr_data_valid = io_data_1_in_26_bits_valid; // @[pe.scala 313:27]
  assign MemController_48_io_wr_data_bits = io_data_1_in_26_bits_bits; // @[pe.scala 313:27]
  assign MemController_49_clock = clock;
  assign MemController_49_reset = reset;
  assign MemController_49_io_rd_valid = io_exec_valid; // @[pe.scala 310:28]
  assign MemController_49_io_wr_valid = io_data_1_in_27_valid; // @[pe.scala 311:28]
  assign MemController_49_io_wr_data_valid = io_data_1_in_27_bits_valid; // @[pe.scala 313:27]
  assign MemController_49_io_wr_data_bits = io_data_1_in_27_bits_bits; // @[pe.scala 313:27]
  assign MemController_50_clock = clock;
  assign MemController_50_reset = reset;
  assign MemController_50_io_rd_valid = io_exec_valid; // @[pe.scala 310:28]
  assign MemController_50_io_wr_valid = io_data_1_in_28_valid; // @[pe.scala 311:28]
  assign MemController_50_io_wr_data_valid = io_data_1_in_28_bits_valid; // @[pe.scala 313:27]
  assign MemController_50_io_wr_data_bits = io_data_1_in_28_bits_bits; // @[pe.scala 313:27]
  assign MemController_51_clock = clock;
  assign MemController_51_reset = reset;
  assign MemController_51_io_rd_valid = io_exec_valid; // @[pe.scala 310:28]
  assign MemController_51_io_wr_valid = io_data_1_in_29_valid; // @[pe.scala 311:28]
  assign MemController_51_io_wr_data_valid = io_data_1_in_29_bits_valid; // @[pe.scala 313:27]
  assign MemController_51_io_wr_data_bits = io_data_1_in_29_bits_bits; // @[pe.scala 313:27]
  assign MemController_52_clock = clock;
  assign MemController_52_reset = reset;
  assign MemController_52_io_rd_valid = io_out_valid; // @[pe.scala 316:28]
  assign MemController_52_io_wr_valid = PENetwork_52_io_to_mem_valid; // @[pe.scala 315:28]
  assign MemController_52_io_wr_data_valid = PENetwork_52_io_to_mem_valid; // @[pe.scala 317:27]
  assign MemController_52_io_wr_data_bits = PENetwork_52_io_to_mem_bits; // @[pe.scala 317:27]
  assign MemController_53_clock = clock;
  assign MemController_53_reset = reset;
  assign MemController_53_io_rd_valid = io_out_valid; // @[pe.scala 316:28]
  assign MemController_53_io_wr_valid = PENetwork_53_io_to_mem_valid; // @[pe.scala 315:28]
  assign MemController_53_io_wr_data_valid = PENetwork_53_io_to_mem_valid; // @[pe.scala 317:27]
  assign MemController_53_io_wr_data_bits = PENetwork_53_io_to_mem_bits; // @[pe.scala 317:27]
  assign MemController_54_clock = clock;
  assign MemController_54_reset = reset;
  assign MemController_54_io_rd_valid = io_out_valid; // @[pe.scala 316:28]
  assign MemController_54_io_wr_valid = PENetwork_54_io_to_mem_valid; // @[pe.scala 315:28]
  assign MemController_54_io_wr_data_valid = PENetwork_54_io_to_mem_valid; // @[pe.scala 317:27]
  assign MemController_54_io_wr_data_bits = PENetwork_54_io_to_mem_bits; // @[pe.scala 317:27]
  assign MemController_55_clock = clock;
  assign MemController_55_reset = reset;
  assign MemController_55_io_rd_valid = io_out_valid; // @[pe.scala 316:28]
  assign MemController_55_io_wr_valid = PENetwork_55_io_to_mem_valid; // @[pe.scala 315:28]
  assign MemController_55_io_wr_data_valid = PENetwork_55_io_to_mem_valid; // @[pe.scala 317:27]
  assign MemController_55_io_wr_data_bits = PENetwork_55_io_to_mem_bits; // @[pe.scala 317:27]
  assign MemController_56_clock = clock;
  assign MemController_56_reset = reset;
  assign MemController_56_io_rd_valid = io_out_valid; // @[pe.scala 316:28]
  assign MemController_56_io_wr_valid = PENetwork_56_io_to_mem_valid; // @[pe.scala 315:28]
  assign MemController_56_io_wr_data_valid = PENetwork_56_io_to_mem_valid; // @[pe.scala 317:27]
  assign MemController_56_io_wr_data_bits = PENetwork_56_io_to_mem_bits; // @[pe.scala 317:27]
  assign MemController_57_clock = clock;
  assign MemController_57_reset = reset;
  assign MemController_57_io_rd_valid = io_out_valid; // @[pe.scala 316:28]
  assign MemController_57_io_wr_valid = PENetwork_57_io_to_mem_valid; // @[pe.scala 315:28]
  assign MemController_57_io_wr_data_valid = PENetwork_57_io_to_mem_valid; // @[pe.scala 317:27]
  assign MemController_57_io_wr_data_bits = PENetwork_57_io_to_mem_bits; // @[pe.scala 317:27]
  assign MemController_58_clock = clock;
  assign MemController_58_reset = reset;
  assign MemController_58_io_rd_valid = io_out_valid; // @[pe.scala 316:28]
  assign MemController_58_io_wr_valid = PENetwork_58_io_to_mem_valid; // @[pe.scala 315:28]
  assign MemController_58_io_wr_data_valid = PENetwork_58_io_to_mem_valid; // @[pe.scala 317:27]
  assign MemController_58_io_wr_data_bits = PENetwork_58_io_to_mem_bits; // @[pe.scala 317:27]
  assign MemController_59_clock = clock;
  assign MemController_59_reset = reset;
  assign MemController_59_io_rd_valid = io_out_valid; // @[pe.scala 316:28]
  assign MemController_59_io_wr_valid = PENetwork_59_io_to_mem_valid; // @[pe.scala 315:28]
  assign MemController_59_io_wr_data_valid = PENetwork_59_io_to_mem_valid; // @[pe.scala 317:27]
  assign MemController_59_io_wr_data_bits = PENetwork_59_io_to_mem_bits; // @[pe.scala 317:27]
  assign MemController_60_clock = clock;
  assign MemController_60_reset = reset;
  assign MemController_60_io_rd_valid = io_out_valid; // @[pe.scala 316:28]
  assign MemController_60_io_wr_valid = PENetwork_60_io_to_mem_valid; // @[pe.scala 315:28]
  assign MemController_60_io_wr_data_valid = PENetwork_60_io_to_mem_valid; // @[pe.scala 317:27]
  assign MemController_60_io_wr_data_bits = PENetwork_60_io_to_mem_bits; // @[pe.scala 317:27]
  assign MemController_61_clock = clock;
  assign MemController_61_reset = reset;
  assign MemController_61_io_rd_valid = io_out_valid; // @[pe.scala 316:28]
  assign MemController_61_io_wr_valid = PENetwork_61_io_to_mem_valid; // @[pe.scala 315:28]
  assign MemController_61_io_wr_data_valid = PENetwork_61_io_to_mem_valid; // @[pe.scala 317:27]
  assign MemController_61_io_wr_data_bits = PENetwork_61_io_to_mem_bits; // @[pe.scala 317:27]
  assign MemController_62_clock = clock;
  assign MemController_62_reset = reset;
  assign MemController_62_io_rd_valid = io_out_valid; // @[pe.scala 316:28]
  assign MemController_62_io_wr_valid = PENetwork_62_io_to_mem_valid; // @[pe.scala 315:28]
  assign MemController_62_io_wr_data_valid = PENetwork_62_io_to_mem_valid; // @[pe.scala 317:27]
  assign MemController_62_io_wr_data_bits = PENetwork_62_io_to_mem_bits; // @[pe.scala 317:27]
  assign MemController_63_clock = clock;
  assign MemController_63_reset = reset;
  assign MemController_63_io_rd_valid = io_out_valid; // @[pe.scala 316:28]
  assign MemController_63_io_wr_valid = PENetwork_63_io_to_mem_valid; // @[pe.scala 315:28]
  assign MemController_63_io_wr_data_valid = PENetwork_63_io_to_mem_valid; // @[pe.scala 317:27]
  assign MemController_63_io_wr_data_bits = PENetwork_63_io_to_mem_bits; // @[pe.scala 317:27]
  assign MemController_64_clock = clock;
  assign MemController_64_reset = reset;
  assign MemController_64_io_rd_valid = io_out_valid; // @[pe.scala 316:28]
  assign MemController_64_io_wr_valid = PENetwork_64_io_to_mem_valid; // @[pe.scala 315:28]
  assign MemController_64_io_wr_data_valid = PENetwork_64_io_to_mem_valid; // @[pe.scala 317:27]
  assign MemController_64_io_wr_data_bits = PENetwork_64_io_to_mem_bits; // @[pe.scala 317:27]
  assign MemController_65_clock = clock;
  assign MemController_65_reset = reset;
  assign MemController_65_io_rd_valid = io_out_valid; // @[pe.scala 316:28]
  assign MemController_65_io_wr_valid = PENetwork_65_io_to_mem_valid; // @[pe.scala 315:28]
  assign MemController_65_io_wr_data_valid = PENetwork_65_io_to_mem_valid; // @[pe.scala 317:27]
  assign MemController_65_io_wr_data_bits = PENetwork_65_io_to_mem_bits; // @[pe.scala 317:27]
  assign MemController_66_clock = clock;
  assign MemController_66_reset = reset;
  assign MemController_66_io_rd_valid = io_out_valid; // @[pe.scala 316:28]
  assign MemController_66_io_wr_valid = PENetwork_66_io_to_mem_valid; // @[pe.scala 315:28]
  assign MemController_66_io_wr_data_valid = PENetwork_66_io_to_mem_valid; // @[pe.scala 317:27]
  assign MemController_66_io_wr_data_bits = PENetwork_66_io_to_mem_bits; // @[pe.scala 317:27]
  assign MemController_67_clock = clock;
  assign MemController_67_reset = reset;
  assign MemController_67_io_rd_valid = io_out_valid; // @[pe.scala 316:28]
  assign MemController_67_io_wr_valid = PENetwork_67_io_to_mem_valid; // @[pe.scala 315:28]
  assign MemController_67_io_wr_data_valid = PENetwork_67_io_to_mem_valid; // @[pe.scala 317:27]
  assign MemController_67_io_wr_data_bits = PENetwork_67_io_to_mem_bits; // @[pe.scala 317:27]
  assign MemController_68_clock = clock;
  assign MemController_68_reset = reset;
  assign MemController_68_io_rd_valid = io_out_valid; // @[pe.scala 316:28]
  assign MemController_68_io_wr_valid = PENetwork_68_io_to_mem_valid; // @[pe.scala 315:28]
  assign MemController_68_io_wr_data_valid = PENetwork_68_io_to_mem_valid; // @[pe.scala 317:27]
  assign MemController_68_io_wr_data_bits = PENetwork_68_io_to_mem_bits; // @[pe.scala 317:27]
  assign MemController_69_clock = clock;
  assign MemController_69_reset = reset;
  assign MemController_69_io_rd_valid = io_out_valid; // @[pe.scala 316:28]
  assign MemController_69_io_wr_valid = PENetwork_69_io_to_mem_valid; // @[pe.scala 315:28]
  assign MemController_69_io_wr_data_valid = PENetwork_69_io_to_mem_valid; // @[pe.scala 317:27]
  assign MemController_69_io_wr_data_bits = PENetwork_69_io_to_mem_bits; // @[pe.scala 317:27]
  assign MemController_70_clock = clock;
  assign MemController_70_reset = reset;
  assign MemController_70_io_rd_valid = io_out_valid; // @[pe.scala 316:28]
  assign MemController_70_io_wr_valid = PENetwork_70_io_to_mem_valid; // @[pe.scala 315:28]
  assign MemController_70_io_wr_data_valid = PENetwork_70_io_to_mem_valid; // @[pe.scala 317:27]
  assign MemController_70_io_wr_data_bits = PENetwork_70_io_to_mem_bits; // @[pe.scala 317:27]
  assign MemController_71_clock = clock;
  assign MemController_71_reset = reset;
  assign MemController_71_io_rd_valid = io_out_valid; // @[pe.scala 316:28]
  assign MemController_71_io_wr_valid = PENetwork_71_io_to_mem_valid; // @[pe.scala 315:28]
  assign MemController_71_io_wr_data_valid = PENetwork_71_io_to_mem_valid; // @[pe.scala 317:27]
  assign MemController_71_io_wr_data_bits = PENetwork_71_io_to_mem_bits; // @[pe.scala 317:27]
  assign MemController_72_clock = clock;
  assign MemController_72_reset = reset;
  assign MemController_72_io_rd_valid = io_out_valid; // @[pe.scala 316:28]
  assign MemController_72_io_wr_valid = PENetwork_72_io_to_mem_valid; // @[pe.scala 315:28]
  assign MemController_72_io_wr_data_valid = PENetwork_72_io_to_mem_valid; // @[pe.scala 317:27]
  assign MemController_72_io_wr_data_bits = PENetwork_72_io_to_mem_bits; // @[pe.scala 317:27]
  assign MemController_73_clock = clock;
  assign MemController_73_reset = reset;
  assign MemController_73_io_rd_valid = io_out_valid; // @[pe.scala 316:28]
  assign MemController_73_io_wr_valid = PENetwork_73_io_to_mem_valid; // @[pe.scala 315:28]
  assign MemController_73_io_wr_data_valid = PENetwork_73_io_to_mem_valid; // @[pe.scala 317:27]
  assign MemController_73_io_wr_data_bits = PENetwork_73_io_to_mem_bits; // @[pe.scala 317:27]
  assign MemController_74_clock = clock;
  assign MemController_74_reset = reset;
  assign MemController_74_io_rd_valid = io_out_valid; // @[pe.scala 316:28]
  assign MemController_74_io_wr_valid = PENetwork_74_io_to_mem_valid; // @[pe.scala 315:28]
  assign MemController_74_io_wr_data_valid = PENetwork_74_io_to_mem_valid; // @[pe.scala 317:27]
  assign MemController_74_io_wr_data_bits = PENetwork_74_io_to_mem_bits; // @[pe.scala 317:27]
  assign MemController_75_clock = clock;
  assign MemController_75_reset = reset;
  assign MemController_75_io_rd_valid = io_out_valid; // @[pe.scala 316:28]
  assign MemController_75_io_wr_valid = PENetwork_75_io_to_mem_valid; // @[pe.scala 315:28]
  assign MemController_75_io_wr_data_valid = PENetwork_75_io_to_mem_valid; // @[pe.scala 317:27]
  assign MemController_75_io_wr_data_bits = PENetwork_75_io_to_mem_bits; // @[pe.scala 317:27]
  assign MemController_76_clock = clock;
  assign MemController_76_reset = reset;
  assign MemController_76_io_rd_valid = io_out_valid; // @[pe.scala 316:28]
  assign MemController_76_io_wr_valid = PENetwork_76_io_to_mem_valid; // @[pe.scala 315:28]
  assign MemController_76_io_wr_data_valid = PENetwork_76_io_to_mem_valid; // @[pe.scala 317:27]
  assign MemController_76_io_wr_data_bits = PENetwork_76_io_to_mem_bits; // @[pe.scala 317:27]
  assign MemController_77_clock = clock;
  assign MemController_77_reset = reset;
  assign MemController_77_io_rd_valid = io_out_valid; // @[pe.scala 316:28]
  assign MemController_77_io_wr_valid = PENetwork_77_io_to_mem_valid; // @[pe.scala 315:28]
  assign MemController_77_io_wr_data_valid = PENetwork_77_io_to_mem_valid; // @[pe.scala 317:27]
  assign MemController_77_io_wr_data_bits = PENetwork_77_io_to_mem_bits; // @[pe.scala 317:27]
  assign MemController_78_clock = clock;
  assign MemController_78_reset = reset;
  assign MemController_78_io_rd_valid = io_out_valid; // @[pe.scala 316:28]
  assign MemController_78_io_wr_valid = PENetwork_78_io_to_mem_valid; // @[pe.scala 315:28]
  assign MemController_78_io_wr_data_valid = PENetwork_78_io_to_mem_valid; // @[pe.scala 317:27]
  assign MemController_78_io_wr_data_bits = PENetwork_78_io_to_mem_bits; // @[pe.scala 317:27]
  assign MemController_79_clock = clock;
  assign MemController_79_reset = reset;
  assign MemController_79_io_rd_valid = io_out_valid; // @[pe.scala 316:28]
  assign MemController_79_io_wr_valid = PENetwork_79_io_to_mem_valid; // @[pe.scala 315:28]
  assign MemController_79_io_wr_data_valid = PENetwork_79_io_to_mem_valid; // @[pe.scala 317:27]
  assign MemController_79_io_wr_data_bits = PENetwork_79_io_to_mem_bits; // @[pe.scala 317:27]
  assign MemController_80_clock = clock;
  assign MemController_80_reset = reset;
  assign MemController_80_io_rd_valid = io_out_valid; // @[pe.scala 316:28]
  assign MemController_80_io_wr_valid = PENetwork_80_io_to_mem_valid; // @[pe.scala 315:28]
  assign MemController_80_io_wr_data_valid = PENetwork_80_io_to_mem_valid; // @[pe.scala 317:27]
  assign MemController_80_io_wr_data_bits = PENetwork_80_io_to_mem_bits; // @[pe.scala 317:27]
  assign MemController_81_clock = clock;
  assign MemController_81_reset = reset;
  assign MemController_81_io_rd_valid = io_out_valid; // @[pe.scala 316:28]
  assign MemController_81_io_wr_valid = PENetwork_81_io_to_mem_valid; // @[pe.scala 315:28]
  assign MemController_81_io_wr_data_valid = PENetwork_81_io_to_mem_valid; // @[pe.scala 317:27]
  assign MemController_81_io_wr_data_bits = PENetwork_81_io_to_mem_bits; // @[pe.scala 317:27]
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"time_ctrl: %d %d %d\n",MultiDimTime_io_index_0,MultiDimTime_io_index_1,MultiDimTime_io_index_2); // @[pe.scala 166:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
