module MultiDimTime(
  input         clock,
  input         reset,
  input         io_in,
  output [1:0]  io_out_0,
  output [1:0]  io_out_1,
  output [1:0]  io_out_2,
  output [15:0] io_index_0,
  output [15:0] io_index_1,
  output [15:0] io_index_2
);
  reg [15:0] regs_0; // @[mem.scala 67:12]
  reg [31:0] _RAND_0;
  reg [15:0] regs_1; // @[mem.scala 67:12]
  reg [31:0] _RAND_1;
  reg [15:0] regs_2; // @[mem.scala 67:12]
  reg [31:0] _RAND_2;
  wire [15:0] _GEN_10 = {{15'd0}, io_in}; // @[mem.scala 69:42]
  wire [15:0] _T_1 = regs_0 + _GEN_10; // @[mem.scala 69:42]
  wire  back_0 = _T_1 == 16'hc; // @[mem.scala 69:48]
  wire [15:0] _T_3 = regs_1 + _GEN_10; // @[mem.scala 69:42]
  wire  next_1 = _T_3 == 16'h10; // @[mem.scala 69:48]
  wire [15:0] _T_5 = regs_2 + _GEN_10; // @[mem.scala 69:42]
  wire  next_2 = _T_5 == 16'h10; // @[mem.scala 69:48]
  wire  back_1 = back_0 & next_1; // @[mem.scala 71:32]
  wire  back_2 = back_1 & next_2; // @[mem.scala 71:32]
  wire  _GEN_1 = back_0 ? 1'h0 : io_in; // @[mem.scala 90:20]
  wire  _GEN_3 = back_1 ? 1'h0 : 1'h1; // @[mem.scala 79:22]
  wire  _GEN_7 = back_2 ? 1'h0 : 1'h1; // @[mem.scala 79:22]
  assign io_out_0 = {{1'd0}, _GEN_1}; // @[mem.scala 92:19 mem.scala 95:19]
  assign io_out_1 = back_0 ? {{1'd0}, _GEN_3} : 2'h2; // @[mem.scala 81:21 mem.scala 84:21 mem.scala 87:19]
  assign io_out_2 = back_1 ? {{1'd0}, _GEN_7} : 2'h2; // @[mem.scala 81:21 mem.scala 84:21 mem.scala 87:19]
  assign io_index_0 = regs_0; // @[mem.scala 76:17]
  assign io_index_1 = regs_1; // @[mem.scala 76:17]
  assign io_index_2 = regs_2; // @[mem.scala 76:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 16'h0;
    end else if (back_0) begin
      regs_0 <= 16'h0;
    end else begin
      regs_0 <= _T_1;
    end
    if (reset) begin
      regs_1 <= 16'h0;
    end else if (back_0) begin
      if (back_1) begin
        regs_1 <= 16'h0;
      end else begin
        regs_1 <= _T_3;
      end
    end
    if (reset) begin
      regs_2 <= 16'h0;
    end else if (back_1) begin
      if (back_2) begin
        regs_2 <= 16'h0;
      end else begin
        regs_2 <= _T_5;
      end
    end
  end
endmodule
module ComputeCellF(
  input          clock,
  input  [255:0] io_data_2_in_bits,
  output         io_data_2_out_valid,
  output [255:0] io_data_2_out_bits,
  input          io_data_1_in_valid,
  input  [255:0] io_data_1_in_bits,
  input          io_data_0_in_valid,
  input  [31:0]  io_data_0_in_bits
);
  wire  My_fmac_aclk; // @[cell.scala 68:62]
  wire  My_fmac_s_axis_a_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_s_axis_a_tdata; // @[cell.scala 68:62]
  wire  My_fmac_s_axis_b_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_s_axis_b_tdata; // @[cell.scala 68:62]
  wire  My_fmac_s_axis_c_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_s_axis_c_tdata; // @[cell.scala 68:62]
  wire  My_fmac_m_axis_result_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_m_axis_result_tdata; // @[cell.scala 68:62]
  wire  My_fmac_1_aclk; // @[cell.scala 68:62]
  wire  My_fmac_1_s_axis_a_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_1_s_axis_a_tdata; // @[cell.scala 68:62]
  wire  My_fmac_1_s_axis_b_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_1_s_axis_b_tdata; // @[cell.scala 68:62]
  wire  My_fmac_1_s_axis_c_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_1_s_axis_c_tdata; // @[cell.scala 68:62]
  wire  My_fmac_1_m_axis_result_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_1_m_axis_result_tdata; // @[cell.scala 68:62]
  wire  My_fmac_2_aclk; // @[cell.scala 68:62]
  wire  My_fmac_2_s_axis_a_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_2_s_axis_a_tdata; // @[cell.scala 68:62]
  wire  My_fmac_2_s_axis_b_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_2_s_axis_b_tdata; // @[cell.scala 68:62]
  wire  My_fmac_2_s_axis_c_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_2_s_axis_c_tdata; // @[cell.scala 68:62]
  wire  My_fmac_2_m_axis_result_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_2_m_axis_result_tdata; // @[cell.scala 68:62]
  wire  My_fmac_3_aclk; // @[cell.scala 68:62]
  wire  My_fmac_3_s_axis_a_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_3_s_axis_a_tdata; // @[cell.scala 68:62]
  wire  My_fmac_3_s_axis_b_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_3_s_axis_b_tdata; // @[cell.scala 68:62]
  wire  My_fmac_3_s_axis_c_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_3_s_axis_c_tdata; // @[cell.scala 68:62]
  wire  My_fmac_3_m_axis_result_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_3_m_axis_result_tdata; // @[cell.scala 68:62]
  wire  My_fmac_4_aclk; // @[cell.scala 68:62]
  wire  My_fmac_4_s_axis_a_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_4_s_axis_a_tdata; // @[cell.scala 68:62]
  wire  My_fmac_4_s_axis_b_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_4_s_axis_b_tdata; // @[cell.scala 68:62]
  wire  My_fmac_4_s_axis_c_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_4_s_axis_c_tdata; // @[cell.scala 68:62]
  wire  My_fmac_4_m_axis_result_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_4_m_axis_result_tdata; // @[cell.scala 68:62]
  wire  My_fmac_5_aclk; // @[cell.scala 68:62]
  wire  My_fmac_5_s_axis_a_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_5_s_axis_a_tdata; // @[cell.scala 68:62]
  wire  My_fmac_5_s_axis_b_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_5_s_axis_b_tdata; // @[cell.scala 68:62]
  wire  My_fmac_5_s_axis_c_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_5_s_axis_c_tdata; // @[cell.scala 68:62]
  wire  My_fmac_5_m_axis_result_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_5_m_axis_result_tdata; // @[cell.scala 68:62]
  wire  My_fmac_6_aclk; // @[cell.scala 68:62]
  wire  My_fmac_6_s_axis_a_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_6_s_axis_a_tdata; // @[cell.scala 68:62]
  wire  My_fmac_6_s_axis_b_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_6_s_axis_b_tdata; // @[cell.scala 68:62]
  wire  My_fmac_6_s_axis_c_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_6_s_axis_c_tdata; // @[cell.scala 68:62]
  wire  My_fmac_6_m_axis_result_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_6_m_axis_result_tdata; // @[cell.scala 68:62]
  wire  My_fmac_7_aclk; // @[cell.scala 68:62]
  wire  My_fmac_7_s_axis_a_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_7_s_axis_a_tdata; // @[cell.scala 68:62]
  wire  My_fmac_7_s_axis_b_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_7_s_axis_b_tdata; // @[cell.scala 68:62]
  wire  My_fmac_7_s_axis_c_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_7_s_axis_c_tdata; // @[cell.scala 68:62]
  wire  My_fmac_7_m_axis_result_tvalid; // @[cell.scala 68:62]
  wire [31:0] My_fmac_7_m_axis_result_tdata; // @[cell.scala 68:62]
  wire [31:0] vec_c_out_1 = My_fmac_1_m_axis_result_tdata; // @[cell.scala 58:25 cell.scala 88:30]
  wire [31:0] vec_c_out_0 = My_fmac_m_axis_result_tdata; // @[cell.scala 58:25 cell.scala 88:30]
  wire [31:0] vec_c_out_3 = My_fmac_3_m_axis_result_tdata; // @[cell.scala 58:25 cell.scala 88:30]
  wire [31:0] vec_c_out_2 = My_fmac_2_m_axis_result_tdata; // @[cell.scala 58:25 cell.scala 88:30]
  wire [127:0] _T_22 = {vec_c_out_3,vec_c_out_2,vec_c_out_1,vec_c_out_0}; // @[cell.scala 91:38]
  wire [31:0] vec_c_out_5 = My_fmac_5_m_axis_result_tdata; // @[cell.scala 58:25 cell.scala 88:30]
  wire [31:0] vec_c_out_4 = My_fmac_4_m_axis_result_tdata; // @[cell.scala 58:25 cell.scala 88:30]
  wire [31:0] vec_c_out_7 = My_fmac_7_m_axis_result_tdata; // @[cell.scala 58:25 cell.scala 88:30]
  wire [31:0] vec_c_out_6 = My_fmac_6_m_axis_result_tdata; // @[cell.scala 58:25 cell.scala 88:30]
  wire [127:0] _T_25 = {vec_c_out_7,vec_c_out_6,vec_c_out_5,vec_c_out_4}; // @[cell.scala 91:38]
  My_fmac My_fmac ( // @[cell.scala 68:62]
    .aclk(My_fmac_aclk),
    .s_axis_a_tvalid(My_fmac_s_axis_a_tvalid),
    .s_axis_a_tdata(My_fmac_s_axis_a_tdata),
    .s_axis_b_tvalid(My_fmac_s_axis_b_tvalid),
    .s_axis_b_tdata(My_fmac_s_axis_b_tdata),
    .s_axis_c_tvalid(My_fmac_s_axis_c_tvalid),
    .s_axis_c_tdata(My_fmac_s_axis_c_tdata),
    .m_axis_result_tvalid(My_fmac_m_axis_result_tvalid),
    .m_axis_result_tdata(My_fmac_m_axis_result_tdata)
  );
  My_fmac My_fmac_1 ( // @[cell.scala 68:62]
    .aclk(My_fmac_1_aclk),
    .s_axis_a_tvalid(My_fmac_1_s_axis_a_tvalid),
    .s_axis_a_tdata(My_fmac_1_s_axis_a_tdata),
    .s_axis_b_tvalid(My_fmac_1_s_axis_b_tvalid),
    .s_axis_b_tdata(My_fmac_1_s_axis_b_tdata),
    .s_axis_c_tvalid(My_fmac_1_s_axis_c_tvalid),
    .s_axis_c_tdata(My_fmac_1_s_axis_c_tdata),
    .m_axis_result_tvalid(My_fmac_1_m_axis_result_tvalid),
    .m_axis_result_tdata(My_fmac_1_m_axis_result_tdata)
  );
  My_fmac My_fmac_2 ( // @[cell.scala 68:62]
    .aclk(My_fmac_2_aclk),
    .s_axis_a_tvalid(My_fmac_2_s_axis_a_tvalid),
    .s_axis_a_tdata(My_fmac_2_s_axis_a_tdata),
    .s_axis_b_tvalid(My_fmac_2_s_axis_b_tvalid),
    .s_axis_b_tdata(My_fmac_2_s_axis_b_tdata),
    .s_axis_c_tvalid(My_fmac_2_s_axis_c_tvalid),
    .s_axis_c_tdata(My_fmac_2_s_axis_c_tdata),
    .m_axis_result_tvalid(My_fmac_2_m_axis_result_tvalid),
    .m_axis_result_tdata(My_fmac_2_m_axis_result_tdata)
  );
  My_fmac My_fmac_3 ( // @[cell.scala 68:62]
    .aclk(My_fmac_3_aclk),
    .s_axis_a_tvalid(My_fmac_3_s_axis_a_tvalid),
    .s_axis_a_tdata(My_fmac_3_s_axis_a_tdata),
    .s_axis_b_tvalid(My_fmac_3_s_axis_b_tvalid),
    .s_axis_b_tdata(My_fmac_3_s_axis_b_tdata),
    .s_axis_c_tvalid(My_fmac_3_s_axis_c_tvalid),
    .s_axis_c_tdata(My_fmac_3_s_axis_c_tdata),
    .m_axis_result_tvalid(My_fmac_3_m_axis_result_tvalid),
    .m_axis_result_tdata(My_fmac_3_m_axis_result_tdata)
  );
  My_fmac My_fmac_4 ( // @[cell.scala 68:62]
    .aclk(My_fmac_4_aclk),
    .s_axis_a_tvalid(My_fmac_4_s_axis_a_tvalid),
    .s_axis_a_tdata(My_fmac_4_s_axis_a_tdata),
    .s_axis_b_tvalid(My_fmac_4_s_axis_b_tvalid),
    .s_axis_b_tdata(My_fmac_4_s_axis_b_tdata),
    .s_axis_c_tvalid(My_fmac_4_s_axis_c_tvalid),
    .s_axis_c_tdata(My_fmac_4_s_axis_c_tdata),
    .m_axis_result_tvalid(My_fmac_4_m_axis_result_tvalid),
    .m_axis_result_tdata(My_fmac_4_m_axis_result_tdata)
  );
  My_fmac My_fmac_5 ( // @[cell.scala 68:62]
    .aclk(My_fmac_5_aclk),
    .s_axis_a_tvalid(My_fmac_5_s_axis_a_tvalid),
    .s_axis_a_tdata(My_fmac_5_s_axis_a_tdata),
    .s_axis_b_tvalid(My_fmac_5_s_axis_b_tvalid),
    .s_axis_b_tdata(My_fmac_5_s_axis_b_tdata),
    .s_axis_c_tvalid(My_fmac_5_s_axis_c_tvalid),
    .s_axis_c_tdata(My_fmac_5_s_axis_c_tdata),
    .m_axis_result_tvalid(My_fmac_5_m_axis_result_tvalid),
    .m_axis_result_tdata(My_fmac_5_m_axis_result_tdata)
  );
  My_fmac My_fmac_6 ( // @[cell.scala 68:62]
    .aclk(My_fmac_6_aclk),
    .s_axis_a_tvalid(My_fmac_6_s_axis_a_tvalid),
    .s_axis_a_tdata(My_fmac_6_s_axis_a_tdata),
    .s_axis_b_tvalid(My_fmac_6_s_axis_b_tvalid),
    .s_axis_b_tdata(My_fmac_6_s_axis_b_tdata),
    .s_axis_c_tvalid(My_fmac_6_s_axis_c_tvalid),
    .s_axis_c_tdata(My_fmac_6_s_axis_c_tdata),
    .m_axis_result_tvalid(My_fmac_6_m_axis_result_tvalid),
    .m_axis_result_tdata(My_fmac_6_m_axis_result_tdata)
  );
  My_fmac My_fmac_7 ( // @[cell.scala 68:62]
    .aclk(My_fmac_7_aclk),
    .s_axis_a_tvalid(My_fmac_7_s_axis_a_tvalid),
    .s_axis_a_tdata(My_fmac_7_s_axis_a_tdata),
    .s_axis_b_tvalid(My_fmac_7_s_axis_b_tvalid),
    .s_axis_b_tdata(My_fmac_7_s_axis_b_tdata),
    .s_axis_c_tvalid(My_fmac_7_s_axis_c_tvalid),
    .s_axis_c_tdata(My_fmac_7_s_axis_c_tdata),
    .m_axis_result_tvalid(My_fmac_7_m_axis_result_tvalid),
    .m_axis_result_tdata(My_fmac_7_m_axis_result_tdata)
  );
  assign io_data_2_out_valid = My_fmac_m_axis_result_tvalid; // @[cell.scala 94:26]
  assign io_data_2_out_bits = {_T_25,_T_22}; // @[cell.scala 91:25]
  assign My_fmac_aclk = clock; // @[cell.scala 81:31]
  assign My_fmac_s_axis_a_tvalid = io_data_0_in_valid; // @[cell.scala 82:41]
  assign My_fmac_s_axis_a_tdata = io_data_0_in_bits; // @[cell.scala 84:40]
  assign My_fmac_s_axis_b_tvalid = io_data_1_in_valid; // @[cell.scala 83:41]
  assign My_fmac_s_axis_b_tdata = io_data_1_in_bits[31:0]; // @[cell.scala 85:40]
  assign My_fmac_s_axis_c_tvalid = 1'h1; // @[cell.scala 86:41]
  assign My_fmac_s_axis_c_tdata = io_data_2_in_bits[31:0]; // @[cell.scala 87:40]
  assign My_fmac_1_aclk = clock; // @[cell.scala 81:31]
  assign My_fmac_1_s_axis_a_tvalid = io_data_0_in_valid; // @[cell.scala 82:41]
  assign My_fmac_1_s_axis_a_tdata = io_data_0_in_bits; // @[cell.scala 84:40]
  assign My_fmac_1_s_axis_b_tvalid = io_data_1_in_valid; // @[cell.scala 83:41]
  assign My_fmac_1_s_axis_b_tdata = io_data_1_in_bits[63:32]; // @[cell.scala 85:40]
  assign My_fmac_1_s_axis_c_tvalid = 1'h1; // @[cell.scala 86:41]
  assign My_fmac_1_s_axis_c_tdata = io_data_2_in_bits[63:32]; // @[cell.scala 87:40]
  assign My_fmac_2_aclk = clock; // @[cell.scala 81:31]
  assign My_fmac_2_s_axis_a_tvalid = io_data_0_in_valid; // @[cell.scala 82:41]
  assign My_fmac_2_s_axis_a_tdata = io_data_0_in_bits; // @[cell.scala 84:40]
  assign My_fmac_2_s_axis_b_tvalid = io_data_1_in_valid; // @[cell.scala 83:41]
  assign My_fmac_2_s_axis_b_tdata = io_data_1_in_bits[95:64]; // @[cell.scala 85:40]
  assign My_fmac_2_s_axis_c_tvalid = 1'h1; // @[cell.scala 86:41]
  assign My_fmac_2_s_axis_c_tdata = io_data_2_in_bits[95:64]; // @[cell.scala 87:40]
  assign My_fmac_3_aclk = clock; // @[cell.scala 81:31]
  assign My_fmac_3_s_axis_a_tvalid = io_data_0_in_valid; // @[cell.scala 82:41]
  assign My_fmac_3_s_axis_a_tdata = io_data_0_in_bits; // @[cell.scala 84:40]
  assign My_fmac_3_s_axis_b_tvalid = io_data_1_in_valid; // @[cell.scala 83:41]
  assign My_fmac_3_s_axis_b_tdata = io_data_1_in_bits[127:96]; // @[cell.scala 85:40]
  assign My_fmac_3_s_axis_c_tvalid = 1'h1; // @[cell.scala 86:41]
  assign My_fmac_3_s_axis_c_tdata = io_data_2_in_bits[127:96]; // @[cell.scala 87:40]
  assign My_fmac_4_aclk = clock; // @[cell.scala 81:31]
  assign My_fmac_4_s_axis_a_tvalid = io_data_0_in_valid; // @[cell.scala 82:41]
  assign My_fmac_4_s_axis_a_tdata = io_data_0_in_bits; // @[cell.scala 84:40]
  assign My_fmac_4_s_axis_b_tvalid = io_data_1_in_valid; // @[cell.scala 83:41]
  assign My_fmac_4_s_axis_b_tdata = io_data_1_in_bits[159:128]; // @[cell.scala 85:40]
  assign My_fmac_4_s_axis_c_tvalid = 1'h1; // @[cell.scala 86:41]
  assign My_fmac_4_s_axis_c_tdata = io_data_2_in_bits[159:128]; // @[cell.scala 87:40]
  assign My_fmac_5_aclk = clock; // @[cell.scala 81:31]
  assign My_fmac_5_s_axis_a_tvalid = io_data_0_in_valid; // @[cell.scala 82:41]
  assign My_fmac_5_s_axis_a_tdata = io_data_0_in_bits; // @[cell.scala 84:40]
  assign My_fmac_5_s_axis_b_tvalid = io_data_1_in_valid; // @[cell.scala 83:41]
  assign My_fmac_5_s_axis_b_tdata = io_data_1_in_bits[191:160]; // @[cell.scala 85:40]
  assign My_fmac_5_s_axis_c_tvalid = 1'h1; // @[cell.scala 86:41]
  assign My_fmac_5_s_axis_c_tdata = io_data_2_in_bits[191:160]; // @[cell.scala 87:40]
  assign My_fmac_6_aclk = clock; // @[cell.scala 81:31]
  assign My_fmac_6_s_axis_a_tvalid = io_data_0_in_valid; // @[cell.scala 82:41]
  assign My_fmac_6_s_axis_a_tdata = io_data_0_in_bits; // @[cell.scala 84:40]
  assign My_fmac_6_s_axis_b_tvalid = io_data_1_in_valid; // @[cell.scala 83:41]
  assign My_fmac_6_s_axis_b_tdata = io_data_1_in_bits[223:192]; // @[cell.scala 85:40]
  assign My_fmac_6_s_axis_c_tvalid = 1'h1; // @[cell.scala 86:41]
  assign My_fmac_6_s_axis_c_tdata = io_data_2_in_bits[223:192]; // @[cell.scala 87:40]
  assign My_fmac_7_aclk = clock; // @[cell.scala 81:31]
  assign My_fmac_7_s_axis_a_tvalid = io_data_0_in_valid; // @[cell.scala 82:41]
  assign My_fmac_7_s_axis_a_tdata = io_data_0_in_bits; // @[cell.scala 84:40]
  assign My_fmac_7_s_axis_b_tvalid = io_data_1_in_valid; // @[cell.scala 83:41]
  assign My_fmac_7_s_axis_b_tdata = io_data_1_in_bits[255:224]; // @[cell.scala 85:40]
  assign My_fmac_7_s_axis_c_tvalid = 1'h1; // @[cell.scala 86:41]
  assign My_fmac_7_s_axis_c_tdata = io_data_2_in_bits[255:224]; // @[cell.scala 87:40]
endmodule
module SystolicInput(
  input         clock,
  input         reset,
  input         io_port_in_valid,
  input  [31:0] io_port_in_bits,
  output        io_port_out_valid,
  output [31:0] io_port_out_bits,
  output        io_to_cell_valid,
  output [31:0] io_to_cell_bits
);
  reg [31:0] reg_bits; // @[pe_modules.scala 55:18]
  reg [31:0] _RAND_0;
  reg  reg_valid; // @[pe_modules.scala 55:18]
  reg [31:0] _RAND_1;
  reg [31:0] to_cell_delay1_bits; // @[pe_modules.scala 55:18]
  reg [31:0] _RAND_2;
  reg  to_cell_delay1_valid; // @[pe_modules.scala 55:18]
  reg [31:0] _RAND_3;
  reg [31:0] to_cell_delay2_bits; // @[pe_modules.scala 55:18]
  reg [31:0] _RAND_4;
  reg  to_cell_delay2_valid; // @[pe_modules.scala 55:18]
  reg [31:0] _RAND_5;
  assign io_port_out_valid = reg_valid; // @[pe_modules.scala 87:15]
  assign io_port_out_bits = reg_bits; // @[pe_modules.scala 87:15]
  assign io_to_cell_valid = to_cell_delay2_valid; // @[pe_modules.scala 88:14]
  assign io_to_cell_bits = to_cell_delay2_bits; // @[pe_modules.scala 88:14]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_bits = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  reg_valid = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  to_cell_delay1_bits = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  to_cell_delay1_valid = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  to_cell_delay2_bits = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  to_cell_delay2_valid = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      reg_bits <= 32'h0;
    end else begin
      reg_bits <= io_port_in_bits;
    end
    if (reset) begin
      reg_valid <= 1'h0;
    end else begin
      reg_valid <= io_port_in_valid;
    end
    if (reset) begin
      to_cell_delay1_bits <= 32'h0;
    end else begin
      to_cell_delay1_bits <= reg_bits;
    end
    if (reset) begin
      to_cell_delay1_valid <= 1'h0;
    end else begin
      to_cell_delay1_valid <= reg_valid;
    end
    if (reset) begin
      to_cell_delay2_bits <= 32'h0;
    end else begin
      to_cell_delay2_bits <= to_cell_delay1_bits;
    end
    if (reset) begin
      to_cell_delay2_valid <= 1'h0;
    end else begin
      to_cell_delay2_valid <= to_cell_delay1_valid;
    end
  end
endmodule
module SystolicInput_1(
  input          clock,
  input          reset,
  input          io_port_in_valid,
  input  [255:0] io_port_in_bits,
  output         io_port_out_valid,
  output [255:0] io_port_out_bits,
  output         io_to_cell_valid,
  output [255:0] io_to_cell_bits
);
  reg [255:0] reg_bits; // @[pe_modules.scala 55:18]
  reg [255:0] _RAND_0;
  reg  reg_valid; // @[pe_modules.scala 55:18]
  reg [31:0] _RAND_1;
  reg [255:0] to_cell_delay1_bits; // @[pe_modules.scala 55:18]
  reg [255:0] _RAND_2;
  reg  to_cell_delay1_valid; // @[pe_modules.scala 55:18]
  reg [31:0] _RAND_3;
  reg [255:0] to_cell_delay2_bits; // @[pe_modules.scala 55:18]
  reg [255:0] _RAND_4;
  reg  to_cell_delay2_valid; // @[pe_modules.scala 55:18]
  reg [31:0] _RAND_5;
  assign io_port_out_valid = reg_valid; // @[pe_modules.scala 87:15]
  assign io_port_out_bits = reg_bits; // @[pe_modules.scala 87:15]
  assign io_to_cell_valid = to_cell_delay2_valid; // @[pe_modules.scala 88:14]
  assign io_to_cell_bits = to_cell_delay2_bits; // @[pe_modules.scala 88:14]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {8{`RANDOM}};
  reg_bits = _RAND_0[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  reg_valid = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {8{`RANDOM}};
  to_cell_delay1_bits = _RAND_2[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  to_cell_delay1_valid = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {8{`RANDOM}};
  to_cell_delay2_bits = _RAND_4[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  to_cell_delay2_valid = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      reg_bits <= 256'h0;
    end else begin
      reg_bits <= io_port_in_bits;
    end
    if (reset) begin
      reg_valid <= 1'h0;
    end else begin
      reg_valid <= io_port_in_valid;
    end
    if (reset) begin
      to_cell_delay1_bits <= 256'h0;
    end else begin
      to_cell_delay1_bits <= reg_bits;
    end
    if (reset) begin
      to_cell_delay1_valid <= 1'h0;
    end else begin
      to_cell_delay1_valid <= reg_valid;
    end
    if (reset) begin
      to_cell_delay2_bits <= 256'h0;
    end else begin
      to_cell_delay2_bits <= to_cell_delay1_bits;
    end
    if (reset) begin
      to_cell_delay2_valid <= 1'h0;
    end else begin
      to_cell_delay2_valid <= to_cell_delay1_valid;
    end
  end
endmodule
module StationaryOutput_InCell(
  input          clock,
  input          reset,
  input          io_port_in_valid,
  input  [255:0] io_port_in_bits,
  output         io_port_out_valid,
  output [255:0] io_port_out_bits,
  input          io_port_sig_stat2trans,
  output         io_port_in_ready,
  input          io_port_out_ready,
  input          io_from_cell_valid,
  input  [255:0] io_from_cell_bits,
  output [255:0] io_to_cell_bits
);
  reg [255:0] trans [0:11]; // @[pe_modules.scala 178:26]
  reg [255:0] _RAND_0;
  wire [255:0] trans_trans_read_data; // @[pe_modules.scala 178:26]
  wire [3:0] trans_trans_read_addr; // @[pe_modules.scala 178:26]
  reg [255:0] _RAND_1;
  wire [255:0] trans__T_3_data; // @[pe_modules.scala 178:26]
  wire [3:0] trans__T_3_addr; // @[pe_modules.scala 178:26]
  wire  trans__T_3_mask; // @[pe_modules.scala 178:26]
  wire  trans__T_3_en; // @[pe_modules.scala 178:26]
  reg  trans_trans_read_en_pipe_0;
  reg [31:0] _RAND_2;
  reg [3:0] trans_trans_read_addr_pipe_0;
  reg [31:0] _RAND_3;
  reg  move_valid; // @[pe_modules.scala 179:21]
  reg [31:0] _RAND_4;
  reg [255:0] move_bits; // @[pe_modules.scala 179:21]
  reg [255:0] _RAND_5;
  reg [255:0] trans_in_addr; // @[pe_modules.scala 180:30]
  reg [255:0] _RAND_6;
  reg [255:0] trans_out_addr; // @[pe_modules.scala 181:31]
  reg [255:0] _RAND_7;
  reg  trans_out_valid; // @[pe_modules.scala 183:32]
  reg [31:0] _RAND_8;
  reg  reg_stat2trans; // @[pe_modules.scala 184:31]
  reg [31:0] _RAND_9;
  wire  _T_1 = reg_stat2trans & io_from_cell_valid; // @[pe_modules.scala 187:22]
  wire  _T_4 = trans_in_addr == 256'hb; // @[pe_modules.scala 189:39]
  wire [255:0] _T_6 = trans_in_addr + 256'h1; // @[pe_modules.scala 189:81]
  wire  _GEN_0 = _T_4 | trans_out_valid; // @[pe_modules.scala 190:47]
  wire  _T_10 = io_port_out_ready & trans_out_valid; // @[pe_modules.scala 198:30]
  wire  _T_11 = trans_out_addr == 256'hb; // @[pe_modules.scala 199:41]
  wire [255:0] _T_13 = trans_out_addr + 256'h1; // @[pe_modules.scala 199:84]
  reg  _T_17; // @[pe_modules.scala 204:15]
  reg [31:0] _RAND_10;
  wire  _GEN_14 = _T_17 | io_port_in_valid; // @[pe_modules.scala 204:58]
  reg  _T_19; // @[pe_modules.scala 210:34]
  reg [31:0] _RAND_11;
  wire  _T_22 = ~reset; // @[pe_modules.scala 214:9]
  assign trans_trans_read_addr = trans_trans_read_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign trans_trans_read_data = trans[trans_trans_read_addr]; // @[pe_modules.scala 178:26]
  `else
  assign trans_trans_read_data = trans_trans_read_addr >= 4'hc ? _RAND_1[255:0] : trans[trans_trans_read_addr]; // @[pe_modules.scala 178:26]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign trans__T_3_data = io_from_cell_bits;
  assign trans__T_3_addr = trans_in_addr[3:0];
  assign trans__T_3_mask = 1'h1;
  assign trans__T_3_en = reg_stat2trans & io_from_cell_valid;
  assign io_port_out_valid = move_valid; // @[pe_modules.scala 211:15]
  assign io_port_out_bits = move_bits; // @[pe_modules.scala 211:15]
  assign io_port_in_ready = _T_19; // @[pe_modules.scala 210:24]
  assign io_to_cell_bits = reg_stat2trans ? 256'h0 : io_from_cell_bits; // @[pe_modules.scala 213:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {8{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 12; initvar = initvar+1)
    trans[initvar] = _RAND_0[255:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {8{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  trans_trans_read_en_pipe_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  trans_trans_read_addr_pipe_0 = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  move_valid = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {8{`RANDOM}};
  move_bits = _RAND_5[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {8{`RANDOM}};
  trans_in_addr = _RAND_6[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {8{`RANDOM}};
  trans_out_addr = _RAND_7[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  trans_out_valid = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  reg_stat2trans = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_17 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_19 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(trans__T_3_en & trans__T_3_mask) begin
      trans[trans__T_3_addr] <= trans__T_3_data; // @[pe_modules.scala 178:26]
    end
    trans_trans_read_en_pipe_0 <= 1'h1;
    trans_trans_read_addr_pipe_0 <= trans_out_addr[3:0];
    if (reset) begin
      move_valid <= 1'h0;
    end else begin
      move_valid <= _GEN_14;
    end
    if (reset) begin
      move_bits <= 256'h0;
    end else if (_T_17) begin
      move_bits <= trans_trans_read_data;
    end else begin
      move_bits <= io_port_in_bits;
    end
    if (reset) begin
      trans_in_addr <= 256'h0;
    end else if (_T_1) begin
      if (_T_4) begin
        trans_in_addr <= 256'h0;
      end else begin
        trans_in_addr <= _T_6;
      end
    end
    if (reset) begin
      trans_out_addr <= 256'h0;
    end else if (_T_10) begin
      if (_T_11) begin
        trans_out_addr <= 256'h0;
      end else begin
        trans_out_addr <= _T_13;
      end
    end
    if (reset) begin
      trans_out_valid <= 1'h0;
    end else if (_T_10) begin
      if (_T_11) begin
        trans_out_valid <= 1'h0;
      end else if (_T_1) begin
        trans_out_valid <= _GEN_0;
      end
    end else if (_T_1) begin
      trans_out_valid <= _GEN_0;
    end
    if (reset) begin
      reg_stat2trans <= 1'h0;
    end else begin
      reg_stat2trans <= io_port_sig_stat2trans;
    end
    _T_17 <= io_port_out_ready & trans_out_valid;
    _T_19 <= ~trans_out_valid;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_22) begin
          $fwrite(32'h80000002,"trans_read: %d, io.port.out_ready.get: %d,trans_out_valid: %d, move: %d %d, pe network out:%d %d\n",trans_trans_read_data,io_port_out_ready,trans_out_valid,move_valid,move_bits,io_port_out_valid,io_port_out_bits); // @[pe_modules.scala 214:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module PE(
  input          clock,
  input          reset,
  input          io_data_2_in_valid,
  input  [255:0] io_data_2_in_bits,
  output         io_data_2_out_valid,
  output [255:0] io_data_2_out_bits,
  input          io_data_2_sig_stat2trans,
  output         io_data_2_in_ready,
  input          io_data_2_out_ready,
  input          io_data_1_in_valid,
  input  [255:0] io_data_1_in_bits,
  output         io_data_1_out_valid,
  output [255:0] io_data_1_out_bits,
  input          io_data_0_in_valid,
  input  [31:0]  io_data_0_in_bits,
  output         io_data_0_out_valid,
  output [31:0]  io_data_0_out_bits
);
  wire  ComputeCellF_clock; // @[pe.scala 44:11]
  wire [255:0] ComputeCellF_io_data_2_in_bits; // @[pe.scala 44:11]
  wire  ComputeCellF_io_data_2_out_valid; // @[pe.scala 44:11]
  wire [255:0] ComputeCellF_io_data_2_out_bits; // @[pe.scala 44:11]
  wire  ComputeCellF_io_data_1_in_valid; // @[pe.scala 44:11]
  wire [255:0] ComputeCellF_io_data_1_in_bits; // @[pe.scala 44:11]
  wire  ComputeCellF_io_data_0_in_valid; // @[pe.scala 44:11]
  wire [31:0] ComputeCellF_io_data_0_in_bits; // @[pe.scala 44:11]
  wire  SystolicInput_clock; // @[pe.scala 46:11]
  wire  SystolicInput_reset; // @[pe.scala 46:11]
  wire  SystolicInput_io_port_in_valid; // @[pe.scala 46:11]
  wire [31:0] SystolicInput_io_port_in_bits; // @[pe.scala 46:11]
  wire  SystolicInput_io_port_out_valid; // @[pe.scala 46:11]
  wire [31:0] SystolicInput_io_port_out_bits; // @[pe.scala 46:11]
  wire  SystolicInput_io_to_cell_valid; // @[pe.scala 46:11]
  wire [31:0] SystolicInput_io_to_cell_bits; // @[pe.scala 46:11]
  wire  SystolicInput_1_clock; // @[pe.scala 46:11]
  wire  SystolicInput_1_reset; // @[pe.scala 46:11]
  wire  SystolicInput_1_io_port_in_valid; // @[pe.scala 46:11]
  wire [255:0] SystolicInput_1_io_port_in_bits; // @[pe.scala 46:11]
  wire  SystolicInput_1_io_port_out_valid; // @[pe.scala 46:11]
  wire [255:0] SystolicInput_1_io_port_out_bits; // @[pe.scala 46:11]
  wire  SystolicInput_1_io_to_cell_valid; // @[pe.scala 46:11]
  wire [255:0] SystolicInput_1_io_to_cell_bits; // @[pe.scala 46:11]
  wire  StationaryOutput_InCell_clock; // @[pe.scala 46:11]
  wire  StationaryOutput_InCell_reset; // @[pe.scala 46:11]
  wire  StationaryOutput_InCell_io_port_in_valid; // @[pe.scala 46:11]
  wire [255:0] StationaryOutput_InCell_io_port_in_bits; // @[pe.scala 46:11]
  wire  StationaryOutput_InCell_io_port_out_valid; // @[pe.scala 46:11]
  wire [255:0] StationaryOutput_InCell_io_port_out_bits; // @[pe.scala 46:11]
  wire  StationaryOutput_InCell_io_port_sig_stat2trans; // @[pe.scala 46:11]
  wire  StationaryOutput_InCell_io_port_in_ready; // @[pe.scala 46:11]
  wire  StationaryOutput_InCell_io_port_out_ready; // @[pe.scala 46:11]
  wire  StationaryOutput_InCell_io_from_cell_valid; // @[pe.scala 46:11]
  wire [255:0] StationaryOutput_InCell_io_from_cell_bits; // @[pe.scala 46:11]
  wire [255:0] StationaryOutput_InCell_io_to_cell_bits; // @[pe.scala 46:11]
  wire  _T_4 = ~reset; // @[pe.scala 56:13]
  ComputeCellF ComputeCellF ( // @[pe.scala 44:11]
    .clock(ComputeCellF_clock),
    .io_data_2_in_bits(ComputeCellF_io_data_2_in_bits),
    .io_data_2_out_valid(ComputeCellF_io_data_2_out_valid),
    .io_data_2_out_bits(ComputeCellF_io_data_2_out_bits),
    .io_data_1_in_valid(ComputeCellF_io_data_1_in_valid),
    .io_data_1_in_bits(ComputeCellF_io_data_1_in_bits),
    .io_data_0_in_valid(ComputeCellF_io_data_0_in_valid),
    .io_data_0_in_bits(ComputeCellF_io_data_0_in_bits)
  );
  SystolicInput SystolicInput ( // @[pe.scala 46:11]
    .clock(SystolicInput_clock),
    .reset(SystolicInput_reset),
    .io_port_in_valid(SystolicInput_io_port_in_valid),
    .io_port_in_bits(SystolicInput_io_port_in_bits),
    .io_port_out_valid(SystolicInput_io_port_out_valid),
    .io_port_out_bits(SystolicInput_io_port_out_bits),
    .io_to_cell_valid(SystolicInput_io_to_cell_valid),
    .io_to_cell_bits(SystolicInput_io_to_cell_bits)
  );
  SystolicInput_1 SystolicInput_1 ( // @[pe.scala 46:11]
    .clock(SystolicInput_1_clock),
    .reset(SystolicInput_1_reset),
    .io_port_in_valid(SystolicInput_1_io_port_in_valid),
    .io_port_in_bits(SystolicInput_1_io_port_in_bits),
    .io_port_out_valid(SystolicInput_1_io_port_out_valid),
    .io_port_out_bits(SystolicInput_1_io_port_out_bits),
    .io_to_cell_valid(SystolicInput_1_io_to_cell_valid),
    .io_to_cell_bits(SystolicInput_1_io_to_cell_bits)
  );
  StationaryOutput_InCell StationaryOutput_InCell ( // @[pe.scala 46:11]
    .clock(StationaryOutput_InCell_clock),
    .reset(StationaryOutput_InCell_reset),
    .io_port_in_valid(StationaryOutput_InCell_io_port_in_valid),
    .io_port_in_bits(StationaryOutput_InCell_io_port_in_bits),
    .io_port_out_valid(StationaryOutput_InCell_io_port_out_valid),
    .io_port_out_bits(StationaryOutput_InCell_io_port_out_bits),
    .io_port_sig_stat2trans(StationaryOutput_InCell_io_port_sig_stat2trans),
    .io_port_in_ready(StationaryOutput_InCell_io_port_in_ready),
    .io_port_out_ready(StationaryOutput_InCell_io_port_out_ready),
    .io_from_cell_valid(StationaryOutput_InCell_io_from_cell_valid),
    .io_from_cell_bits(StationaryOutput_InCell_io_from_cell_bits),
    .io_to_cell_bits(StationaryOutput_InCell_io_to_cell_bits)
  );
  assign io_data_2_out_valid = StationaryOutput_InCell_io_port_out_valid; // @[pe.scala 51:17]
  assign io_data_2_out_bits = StationaryOutput_InCell_io_port_out_bits; // @[pe.scala 51:17]
  assign io_data_2_in_ready = StationaryOutput_InCell_io_port_in_ready; // @[pe.scala 51:17]
  assign io_data_1_out_valid = SystolicInput_1_io_port_out_valid; // @[pe.scala 51:17]
  assign io_data_1_out_bits = SystolicInput_1_io_port_out_bits; // @[pe.scala 51:17]
  assign io_data_0_out_valid = SystolicInput_io_port_out_valid; // @[pe.scala 51:17]
  assign io_data_0_out_bits = SystolicInput_io_port_out_bits; // @[pe.scala 51:17]
  assign ComputeCellF_clock = clock;
  assign ComputeCellF_io_data_2_in_bits = StationaryOutput_InCell_io_to_cell_bits; // @[pe.scala 52:19]
  assign ComputeCellF_io_data_1_in_valid = SystolicInput_1_io_to_cell_valid; // @[pe.scala 52:19]
  assign ComputeCellF_io_data_1_in_bits = SystolicInput_1_io_to_cell_bits; // @[pe.scala 52:19]
  assign ComputeCellF_io_data_0_in_valid = SystolicInput_io_to_cell_valid; // @[pe.scala 52:19]
  assign ComputeCellF_io_data_0_in_bits = SystolicInput_io_to_cell_bits; // @[pe.scala 52:19]
  assign SystolicInput_clock = clock;
  assign SystolicInput_reset = reset;
  assign SystolicInput_io_port_in_valid = io_data_0_in_valid; // @[pe.scala 51:17]
  assign SystolicInput_io_port_in_bits = io_data_0_in_bits; // @[pe.scala 51:17]
  assign SystolicInput_1_clock = clock;
  assign SystolicInput_1_reset = reset;
  assign SystolicInput_1_io_port_in_valid = io_data_1_in_valid; // @[pe.scala 51:17]
  assign SystolicInput_1_io_port_in_bits = io_data_1_in_bits; // @[pe.scala 51:17]
  assign StationaryOutput_InCell_clock = clock;
  assign StationaryOutput_InCell_reset = reset;
  assign StationaryOutput_InCell_io_port_in_valid = io_data_2_in_valid; // @[pe.scala 51:17]
  assign StationaryOutput_InCell_io_port_in_bits = io_data_2_in_bits; // @[pe.scala 51:17]
  assign StationaryOutput_InCell_io_port_sig_stat2trans = io_data_2_sig_stat2trans; // @[pe.scala 51:17 pe.scala 61:38]
  assign StationaryOutput_InCell_io_port_out_ready = io_data_2_out_ready; // @[pe.scala 51:17]
  assign StationaryOutput_InCell_io_from_cell_valid = ComputeCellF_io_data_2_out_valid; // @[pe.scala 54:28]
  assign StationaryOutput_InCell_io_from_cell_bits = ComputeCellF_io_data_2_out_bits; // @[pe.scala 54:28]
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_4) begin
          $fwrite(32'h80000002,"pe out:%d %d\n",StationaryOutput_InCell_io_from_cell_bits,StationaryOutput_InCell_io_from_cell_valid); // @[pe.scala 56:13]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module PENetwork(
  output        io_to_pes_0_in_valid,
  output [31:0] io_to_pes_0_in_bits,
  input         io_to_pes_0_out_valid,
  input  [31:0] io_to_pes_0_out_bits,
  output        io_to_pes_1_in_valid,
  output [31:0] io_to_pes_1_in_bits,
  input         io_to_pes_1_out_valid,
  input  [31:0] io_to_pes_1_out_bits,
  output        io_to_pes_2_in_valid,
  output [31:0] io_to_pes_2_in_bits,
  input         io_to_pes_2_out_valid,
  input  [31:0] io_to_pes_2_out_bits,
  output        io_to_pes_3_in_valid,
  output [31:0] io_to_pes_3_in_bits,
  input         io_to_pes_3_out_valid,
  input  [31:0] io_to_pes_3_out_bits,
  output        io_to_pes_4_in_valid,
  output [31:0] io_to_pes_4_in_bits,
  input         io_to_pes_4_out_valid,
  input  [31:0] io_to_pes_4_out_bits,
  output        io_to_pes_5_in_valid,
  output [31:0] io_to_pes_5_in_bits,
  input         io_to_pes_5_out_valid,
  input  [31:0] io_to_pes_5_out_bits,
  output        io_to_pes_6_in_valid,
  output [31:0] io_to_pes_6_in_bits,
  input         io_to_pes_6_out_valid,
  input  [31:0] io_to_pes_6_out_bits,
  output        io_to_pes_7_in_valid,
  output [31:0] io_to_pes_7_in_bits,
  input         io_to_pes_7_out_valid,
  input  [31:0] io_to_pes_7_out_bits,
  output        io_to_pes_8_in_valid,
  output [31:0] io_to_pes_8_in_bits,
  input         io_to_pes_8_out_valid,
  input  [31:0] io_to_pes_8_out_bits,
  output        io_to_pes_9_in_valid,
  output [31:0] io_to_pes_9_in_bits,
  input         io_to_pes_9_out_valid,
  input  [31:0] io_to_pes_9_out_bits,
  output        io_to_pes_10_in_valid,
  output [31:0] io_to_pes_10_in_bits,
  input         io_to_pes_10_out_valid,
  input  [31:0] io_to_pes_10_out_bits,
  output        io_to_pes_11_in_valid,
  output [31:0] io_to_pes_11_in_bits,
  input         io_to_pes_11_out_valid,
  input  [31:0] io_to_pes_11_out_bits,
  output        io_to_pes_12_in_valid,
  output [31:0] io_to_pes_12_in_bits,
  input         io_to_pes_12_out_valid,
  input  [31:0] io_to_pes_12_out_bits,
  output        io_to_pes_13_in_valid,
  output [31:0] io_to_pes_13_in_bits,
  input         io_to_pes_13_out_valid,
  input  [31:0] io_to_pes_13_out_bits,
  output        io_to_pes_14_in_valid,
  output [31:0] io_to_pes_14_in_bits,
  input         io_to_mem_valid,
  input  [31:0] io_to_mem_bits
);
  assign io_to_pes_0_in_valid = io_to_mem_valid; // @[pe.scala 125:23]
  assign io_to_pes_0_in_bits = io_to_mem_bits; // @[pe.scala 125:23]
  assign io_to_pes_1_in_valid = io_to_pes_0_out_valid; // @[pe.scala 122:23]
  assign io_to_pes_1_in_bits = io_to_pes_0_out_bits; // @[pe.scala 122:23]
  assign io_to_pes_2_in_valid = io_to_pes_1_out_valid; // @[pe.scala 122:23]
  assign io_to_pes_2_in_bits = io_to_pes_1_out_bits; // @[pe.scala 122:23]
  assign io_to_pes_3_in_valid = io_to_pes_2_out_valid; // @[pe.scala 122:23]
  assign io_to_pes_3_in_bits = io_to_pes_2_out_bits; // @[pe.scala 122:23]
  assign io_to_pes_4_in_valid = io_to_pes_3_out_valid; // @[pe.scala 122:23]
  assign io_to_pes_4_in_bits = io_to_pes_3_out_bits; // @[pe.scala 122:23]
  assign io_to_pes_5_in_valid = io_to_pes_4_out_valid; // @[pe.scala 122:23]
  assign io_to_pes_5_in_bits = io_to_pes_4_out_bits; // @[pe.scala 122:23]
  assign io_to_pes_6_in_valid = io_to_pes_5_out_valid; // @[pe.scala 122:23]
  assign io_to_pes_6_in_bits = io_to_pes_5_out_bits; // @[pe.scala 122:23]
  assign io_to_pes_7_in_valid = io_to_pes_6_out_valid; // @[pe.scala 122:23]
  assign io_to_pes_7_in_bits = io_to_pes_6_out_bits; // @[pe.scala 122:23]
  assign io_to_pes_8_in_valid = io_to_pes_7_out_valid; // @[pe.scala 122:23]
  assign io_to_pes_8_in_bits = io_to_pes_7_out_bits; // @[pe.scala 122:23]
  assign io_to_pes_9_in_valid = io_to_pes_8_out_valid; // @[pe.scala 122:23]
  assign io_to_pes_9_in_bits = io_to_pes_8_out_bits; // @[pe.scala 122:23]
  assign io_to_pes_10_in_valid = io_to_pes_9_out_valid; // @[pe.scala 122:23]
  assign io_to_pes_10_in_bits = io_to_pes_9_out_bits; // @[pe.scala 122:23]
  assign io_to_pes_11_in_valid = io_to_pes_10_out_valid; // @[pe.scala 122:23]
  assign io_to_pes_11_in_bits = io_to_pes_10_out_bits; // @[pe.scala 122:23]
  assign io_to_pes_12_in_valid = io_to_pes_11_out_valid; // @[pe.scala 122:23]
  assign io_to_pes_12_in_bits = io_to_pes_11_out_bits; // @[pe.scala 122:23]
  assign io_to_pes_13_in_valid = io_to_pes_12_out_valid; // @[pe.scala 122:23]
  assign io_to_pes_13_in_bits = io_to_pes_12_out_bits; // @[pe.scala 122:23]
  assign io_to_pes_14_in_valid = io_to_pes_13_out_valid; // @[pe.scala 122:23]
  assign io_to_pes_14_in_bits = io_to_pes_13_out_bits; // @[pe.scala 122:23]
endmodule
module PENetwork_11(
  output         io_to_pes_0_in_valid,
  output [255:0] io_to_pes_0_in_bits,
  input          io_to_pes_0_out_valid,
  input  [255:0] io_to_pes_0_out_bits,
  output         io_to_pes_1_in_valid,
  output [255:0] io_to_pes_1_in_bits,
  input          io_to_pes_1_out_valid,
  input  [255:0] io_to_pes_1_out_bits,
  output         io_to_pes_2_in_valid,
  output [255:0] io_to_pes_2_in_bits,
  input          io_to_pes_2_out_valid,
  input  [255:0] io_to_pes_2_out_bits,
  output         io_to_pes_3_in_valid,
  output [255:0] io_to_pes_3_in_bits,
  input          io_to_pes_3_out_valid,
  input  [255:0] io_to_pes_3_out_bits,
  output         io_to_pes_4_in_valid,
  output [255:0] io_to_pes_4_in_bits,
  input          io_to_pes_4_out_valid,
  input  [255:0] io_to_pes_4_out_bits,
  output         io_to_pes_5_in_valid,
  output [255:0] io_to_pes_5_in_bits,
  input          io_to_pes_5_out_valid,
  input  [255:0] io_to_pes_5_out_bits,
  output         io_to_pes_6_in_valid,
  output [255:0] io_to_pes_6_in_bits,
  input          io_to_pes_6_out_valid,
  input  [255:0] io_to_pes_6_out_bits,
  output         io_to_pes_7_in_valid,
  output [255:0] io_to_pes_7_in_bits,
  input          io_to_pes_7_out_valid,
  input  [255:0] io_to_pes_7_out_bits,
  output         io_to_pes_8_in_valid,
  output [255:0] io_to_pes_8_in_bits,
  input          io_to_pes_8_out_valid,
  input  [255:0] io_to_pes_8_out_bits,
  output         io_to_pes_9_in_valid,
  output [255:0] io_to_pes_9_in_bits,
  input          io_to_pes_9_out_valid,
  input  [255:0] io_to_pes_9_out_bits,
  output         io_to_pes_10_in_valid,
  output [255:0] io_to_pes_10_in_bits,
  input          io_to_mem_valid,
  input  [255:0] io_to_mem_bits
);
  assign io_to_pes_0_in_valid = io_to_mem_valid; // @[pe.scala 125:23]
  assign io_to_pes_0_in_bits = io_to_mem_bits; // @[pe.scala 125:23]
  assign io_to_pes_1_in_valid = io_to_pes_0_out_valid; // @[pe.scala 122:23]
  assign io_to_pes_1_in_bits = io_to_pes_0_out_bits; // @[pe.scala 122:23]
  assign io_to_pes_2_in_valid = io_to_pes_1_out_valid; // @[pe.scala 122:23]
  assign io_to_pes_2_in_bits = io_to_pes_1_out_bits; // @[pe.scala 122:23]
  assign io_to_pes_3_in_valid = io_to_pes_2_out_valid; // @[pe.scala 122:23]
  assign io_to_pes_3_in_bits = io_to_pes_2_out_bits; // @[pe.scala 122:23]
  assign io_to_pes_4_in_valid = io_to_pes_3_out_valid; // @[pe.scala 122:23]
  assign io_to_pes_4_in_bits = io_to_pes_3_out_bits; // @[pe.scala 122:23]
  assign io_to_pes_5_in_valid = io_to_pes_4_out_valid; // @[pe.scala 122:23]
  assign io_to_pes_5_in_bits = io_to_pes_4_out_bits; // @[pe.scala 122:23]
  assign io_to_pes_6_in_valid = io_to_pes_5_out_valid; // @[pe.scala 122:23]
  assign io_to_pes_6_in_bits = io_to_pes_5_out_bits; // @[pe.scala 122:23]
  assign io_to_pes_7_in_valid = io_to_pes_6_out_valid; // @[pe.scala 122:23]
  assign io_to_pes_7_in_bits = io_to_pes_6_out_bits; // @[pe.scala 122:23]
  assign io_to_pes_8_in_valid = io_to_pes_7_out_valid; // @[pe.scala 122:23]
  assign io_to_pes_8_in_bits = io_to_pes_7_out_bits; // @[pe.scala 122:23]
  assign io_to_pes_9_in_valid = io_to_pes_8_out_valid; // @[pe.scala 122:23]
  assign io_to_pes_9_in_bits = io_to_pes_8_out_bits; // @[pe.scala 122:23]
  assign io_to_pes_10_in_valid = io_to_pes_9_out_valid; // @[pe.scala 122:23]
  assign io_to_pes_10_in_bits = io_to_pes_9_out_bits; // @[pe.scala 122:23]
endmodule
module PENetwork_26(
  input          clock,
  input          io_to_pes_0_out_valid,
  input  [255:0] io_to_pes_0_out_bits,
  output         io_to_pes_0_sig_stat2trans,
  output         io_to_pes_0_out_ready,
  output         io_to_pes_1_in_valid,
  output [255:0] io_to_pes_1_in_bits,
  input          io_to_pes_1_out_valid,
  input  [255:0] io_to_pes_1_out_bits,
  output         io_to_pes_1_sig_stat2trans,
  input          io_to_pes_1_in_ready,
  output         io_to_pes_1_out_ready,
  output         io_to_pes_2_in_valid,
  output [255:0] io_to_pes_2_in_bits,
  input          io_to_pes_2_out_valid,
  input  [255:0] io_to_pes_2_out_bits,
  output         io_to_pes_2_sig_stat2trans,
  input          io_to_pes_2_in_ready,
  output         io_to_pes_2_out_ready,
  output         io_to_pes_3_in_valid,
  output [255:0] io_to_pes_3_in_bits,
  input          io_to_pes_3_out_valid,
  input  [255:0] io_to_pes_3_out_bits,
  output         io_to_pes_3_sig_stat2trans,
  input          io_to_pes_3_in_ready,
  output         io_to_pes_3_out_ready,
  output         io_to_pes_4_in_valid,
  output [255:0] io_to_pes_4_in_bits,
  input          io_to_pes_4_out_valid,
  input  [255:0] io_to_pes_4_out_bits,
  output         io_to_pes_4_sig_stat2trans,
  input          io_to_pes_4_in_ready,
  output         io_to_pes_4_out_ready,
  output         io_to_pes_5_in_valid,
  output [255:0] io_to_pes_5_in_bits,
  input          io_to_pes_5_out_valid,
  input  [255:0] io_to_pes_5_out_bits,
  output         io_to_pes_5_sig_stat2trans,
  input          io_to_pes_5_in_ready,
  output         io_to_pes_5_out_ready,
  output         io_to_pes_6_in_valid,
  output [255:0] io_to_pes_6_in_bits,
  input          io_to_pes_6_out_valid,
  input  [255:0] io_to_pes_6_out_bits,
  output         io_to_pes_6_sig_stat2trans,
  input          io_to_pes_6_in_ready,
  output         io_to_pes_6_out_ready,
  output         io_to_pes_7_in_valid,
  output [255:0] io_to_pes_7_in_bits,
  input          io_to_pes_7_out_valid,
  input  [255:0] io_to_pes_7_out_bits,
  output         io_to_pes_7_sig_stat2trans,
  input          io_to_pes_7_in_ready,
  output         io_to_pes_7_out_ready,
  output         io_to_pes_8_in_valid,
  output [255:0] io_to_pes_8_in_bits,
  input          io_to_pes_8_out_valid,
  input  [255:0] io_to_pes_8_out_bits,
  output         io_to_pes_8_sig_stat2trans,
  input          io_to_pes_8_in_ready,
  output         io_to_pes_8_out_ready,
  output         io_to_pes_9_in_valid,
  output [255:0] io_to_pes_9_in_bits,
  input          io_to_pes_9_out_valid,
  input  [255:0] io_to_pes_9_out_bits,
  output         io_to_pes_9_sig_stat2trans,
  input          io_to_pes_9_in_ready,
  output         io_to_pes_9_out_ready,
  output         io_to_pes_10_in_valid,
  output [255:0] io_to_pes_10_in_bits,
  input          io_to_pes_10_out_valid,
  input  [255:0] io_to_pes_10_out_bits,
  output         io_to_pes_10_sig_stat2trans,
  input          io_to_pes_10_in_ready,
  output         io_to_mem_valid,
  output [255:0] io_to_mem_bits,
  input          io_sig_stat2trans
);
  reg  _T; // @[Reg.scala 15:16]
  reg [31:0] _RAND_0;
  reg  _T_1; // @[Reg.scala 15:16]
  reg [31:0] _RAND_1;
  reg  _T_2; // @[Reg.scala 15:16]
  reg [31:0] _RAND_2;
  reg  _T_3; // @[Reg.scala 15:16]
  reg [31:0] _RAND_3;
  reg  _T_4; // @[Reg.scala 15:16]
  reg [31:0] _RAND_4;
  reg  _T_5; // @[Reg.scala 15:16]
  reg [31:0] _RAND_5;
  reg  _T_6; // @[Reg.scala 15:16]
  reg [31:0] _RAND_6;
  reg  _T_7; // @[Reg.scala 15:16]
  reg [31:0] _RAND_7;
  reg  _T_8; // @[Reg.scala 15:16]
  reg [31:0] _RAND_8;
  reg  _T_9; // @[Reg.scala 15:16]
  reg [31:0] _RAND_9;
  reg  _T_10; // @[Reg.scala 15:16]
  reg [31:0] _RAND_10;
  reg  _T_11; // @[Reg.scala 15:16]
  reg [31:0] _RAND_11;
  reg  _T_12; // @[Reg.scala 15:16]
  reg [31:0] _RAND_12;
  reg  _T_13; // @[Reg.scala 15:16]
  reg [31:0] _RAND_13;
  reg  _T_14; // @[Reg.scala 15:16]
  reg [31:0] _RAND_14;
  reg  _T_15; // @[Reg.scala 15:16]
  reg [31:0] _RAND_15;
  reg  _T_16; // @[Reg.scala 15:16]
  reg [31:0] _RAND_16;
  reg  _T_17; // @[Reg.scala 15:16]
  reg [31:0] _RAND_17;
  reg  _T_18; // @[Reg.scala 15:16]
  reg [31:0] _RAND_18;
  reg  _T_19; // @[Reg.scala 15:16]
  reg [31:0] _RAND_19;
  reg  _T_20; // @[Reg.scala 15:16]
  reg [31:0] _RAND_20;
  reg  _T_21; // @[Reg.scala 15:16]
  reg [31:0] _RAND_21;
  reg  _T_22; // @[Reg.scala 15:16]
  reg [31:0] _RAND_22;
  reg  _T_23; // @[Reg.scala 15:16]
  reg [31:0] _RAND_23;
  reg  _T_24; // @[Reg.scala 15:16]
  reg [31:0] _RAND_24;
  reg  _T_25; // @[Reg.scala 15:16]
  reg [31:0] _RAND_25;
  reg  _T_26; // @[Reg.scala 15:16]
  reg [31:0] _RAND_26;
  reg  _T_27; // @[Reg.scala 15:16]
  reg [31:0] _RAND_27;
  reg  _T_28; // @[Reg.scala 15:16]
  reg [31:0] _RAND_28;
  reg  _T_29; // @[Reg.scala 15:16]
  reg [31:0] _RAND_29;
  reg  _T_30; // @[Reg.scala 15:16]
  reg [31:0] _RAND_30;
  reg  _T_31; // @[Reg.scala 15:16]
  reg [31:0] _RAND_31;
  reg  _T_32; // @[Reg.scala 15:16]
  reg [31:0] _RAND_32;
  reg  _T_33; // @[Reg.scala 15:16]
  reg [31:0] _RAND_33;
  reg  _T_34; // @[Reg.scala 15:16]
  reg [31:0] _RAND_34;
  reg  _T_35; // @[Reg.scala 15:16]
  reg [31:0] _RAND_35;
  reg  _T_36; // @[Reg.scala 15:16]
  reg [31:0] _RAND_36;
  reg  _T_37; // @[Reg.scala 15:16]
  reg [31:0] _RAND_37;
  reg  _T_38; // @[Reg.scala 15:16]
  reg [31:0] _RAND_38;
  reg  _T_39; // @[Reg.scala 15:16]
  reg [31:0] _RAND_39;
  reg  _T_40; // @[Reg.scala 15:16]
  reg [31:0] _RAND_40;
  reg  _T_41; // @[Reg.scala 15:16]
  reg [31:0] _RAND_41;
  reg  _T_42; // @[Reg.scala 15:16]
  reg [31:0] _RAND_42;
  reg  _T_43; // @[Reg.scala 15:16]
  reg [31:0] _RAND_43;
  reg  _T_44; // @[Reg.scala 15:16]
  reg [31:0] _RAND_44;
  reg  _T_45; // @[Reg.scala 15:16]
  reg [31:0] _RAND_45;
  reg  _T_46; // @[Reg.scala 15:16]
  reg [31:0] _RAND_46;
  reg  _T_47; // @[Reg.scala 15:16]
  reg [31:0] _RAND_47;
  reg  _T_48; // @[Reg.scala 15:16]
  reg [31:0] _RAND_48;
  reg  _T_49; // @[Reg.scala 15:16]
  reg [31:0] _RAND_49;
  reg  _T_50; // @[Reg.scala 15:16]
  reg [31:0] _RAND_50;
  reg  _T_51; // @[Reg.scala 15:16]
  reg [31:0] _RAND_51;
  reg  _T_52; // @[Reg.scala 15:16]
  reg [31:0] _RAND_52;
  reg  _T_53; // @[Reg.scala 15:16]
  reg [31:0] _RAND_53;
  reg  _T_54; // @[Reg.scala 15:16]
  reg [31:0] _RAND_54;
  reg  _T_55; // @[Reg.scala 15:16]
  reg [31:0] _RAND_55;
  reg  _T_56; // @[Reg.scala 15:16]
  reg [31:0] _RAND_56;
  reg  _T_57; // @[Reg.scala 15:16]
  reg [31:0] _RAND_57;
  reg  _T_58; // @[Reg.scala 15:16]
  reg [31:0] _RAND_58;
  reg  _T_59; // @[Reg.scala 15:16]
  reg [31:0] _RAND_59;
  reg  _T_60; // @[Reg.scala 15:16]
  reg [31:0] _RAND_60;
  reg  _T_61; // @[Reg.scala 15:16]
  reg [31:0] _RAND_61;
  reg  _T_62; // @[Reg.scala 15:16]
  reg [31:0] _RAND_62;
  reg  _T_63; // @[Reg.scala 15:16]
  reg [31:0] _RAND_63;
  reg  _T_64; // @[Reg.scala 15:16]
  reg [31:0] _RAND_64;
  reg  _T_65; // @[Reg.scala 15:16]
  reg [31:0] _RAND_65;
  reg  _T_66; // @[Reg.scala 15:16]
  reg [31:0] _RAND_66;
  reg  _T_67; // @[Reg.scala 15:16]
  reg [31:0] _RAND_67;
  reg  _T_68; // @[Reg.scala 15:16]
  reg [31:0] _RAND_68;
  reg  _T_69; // @[Reg.scala 15:16]
  reg [31:0] _RAND_69;
  reg  _T_70; // @[Reg.scala 15:16]
  reg [31:0] _RAND_70;
  reg  _T_71; // @[Reg.scala 15:16]
  reg [31:0] _RAND_71;
  reg  _T_72; // @[Reg.scala 15:16]
  reg [31:0] _RAND_72;
  reg  _T_73; // @[Reg.scala 15:16]
  reg [31:0] _RAND_73;
  reg  _T_74; // @[Reg.scala 15:16]
  reg [31:0] _RAND_74;
  reg  _T_75; // @[Reg.scala 15:16]
  reg [31:0] _RAND_75;
  reg  _T_76; // @[Reg.scala 15:16]
  reg [31:0] _RAND_76;
  reg  _T_77; // @[Reg.scala 15:16]
  reg [31:0] _RAND_77;
  reg  _T_78; // @[Reg.scala 15:16]
  reg [31:0] _RAND_78;
  reg  _T_79; // @[Reg.scala 15:16]
  reg [31:0] _RAND_79;
  reg  _T_80; // @[Reg.scala 15:16]
  reg [31:0] _RAND_80;
  reg  _T_81; // @[Reg.scala 15:16]
  reg [31:0] _RAND_81;
  reg  _T_82; // @[Reg.scala 15:16]
  reg [31:0] _RAND_82;
  reg  _T_83; // @[Reg.scala 15:16]
  reg [31:0] _RAND_83;
  reg  _T_84; // @[Reg.scala 15:16]
  reg [31:0] _RAND_84;
  reg  _T_85; // @[Reg.scala 15:16]
  reg [31:0] _RAND_85;
  reg  _T_86; // @[Reg.scala 15:16]
  reg [31:0] _RAND_86;
  reg  _T_87; // @[Reg.scala 15:16]
  reg [31:0] _RAND_87;
  reg  _T_88; // @[Reg.scala 15:16]
  reg [31:0] _RAND_88;
  reg  _T_89; // @[Reg.scala 15:16]
  reg [31:0] _RAND_89;
  reg  _T_90; // @[Reg.scala 15:16]
  reg [31:0] _RAND_90;
  reg  _T_91; // @[Reg.scala 15:16]
  reg [31:0] _RAND_91;
  reg  _T_92; // @[Reg.scala 15:16]
  reg [31:0] _RAND_92;
  reg  _T_93; // @[Reg.scala 15:16]
  reg [31:0] _RAND_93;
  reg  _T_94; // @[Reg.scala 15:16]
  reg [31:0] _RAND_94;
  reg  _T_95; // @[Reg.scala 15:16]
  reg [31:0] _RAND_95;
  reg  _T_96; // @[Reg.scala 15:16]
  reg [31:0] _RAND_96;
  reg  _T_97; // @[Reg.scala 15:16]
  reg [31:0] _RAND_97;
  reg  _T_98; // @[Reg.scala 15:16]
  reg [31:0] _RAND_98;
  reg  _T_99; // @[Reg.scala 15:16]
  reg [31:0] _RAND_99;
  reg  _T_100; // @[Reg.scala 15:16]
  reg [31:0] _RAND_100;
  reg  _T_101; // @[Reg.scala 15:16]
  reg [31:0] _RAND_101;
  reg  _T_102; // @[Reg.scala 15:16]
  reg [31:0] _RAND_102;
  reg  _T_103; // @[Reg.scala 15:16]
  reg [31:0] _RAND_103;
  reg  _T_104; // @[Reg.scala 15:16]
  reg [31:0] _RAND_104;
  reg  _T_105; // @[Reg.scala 15:16]
  reg [31:0] _RAND_105;
  reg  _T_106; // @[Reg.scala 15:16]
  reg [31:0] _RAND_106;
  reg  _T_107; // @[Reg.scala 15:16]
  reg [31:0] _RAND_107;
  reg  _T_108; // @[Reg.scala 15:16]
  reg [31:0] _RAND_108;
  reg  _T_109; // @[Reg.scala 15:16]
  reg [31:0] _RAND_109;
  reg  _T_110; // @[Reg.scala 15:16]
  reg [31:0] _RAND_110;
  reg  _T_111; // @[Reg.scala 15:16]
  reg [31:0] _RAND_111;
  reg  _T_112; // @[Reg.scala 15:16]
  reg [31:0] _RAND_112;
  reg  _T_113; // @[Reg.scala 15:16]
  reg [31:0] _RAND_113;
  reg  _T_114; // @[Reg.scala 15:16]
  reg [31:0] _RAND_114;
  reg  _T_115; // @[Reg.scala 15:16]
  reg [31:0] _RAND_115;
  reg  _T_116; // @[Reg.scala 15:16]
  reg [31:0] _RAND_116;
  reg  _T_117; // @[Reg.scala 15:16]
  reg [31:0] _RAND_117;
  reg  _T_118; // @[Reg.scala 15:16]
  reg [31:0] _RAND_118;
  reg  _T_119; // @[Reg.scala 15:16]
  reg [31:0] _RAND_119;
  reg  _T_120; // @[Reg.scala 15:16]
  reg [31:0] _RAND_120;
  reg  _T_121; // @[Reg.scala 15:16]
  reg [31:0] _RAND_121;
  reg  _T_122; // @[Reg.scala 15:16]
  reg [31:0] _RAND_122;
  reg  _T_123; // @[Reg.scala 15:16]
  reg [31:0] _RAND_123;
  reg  _T_124; // @[Reg.scala 15:16]
  reg [31:0] _RAND_124;
  reg  _T_125; // @[Reg.scala 15:16]
  reg [31:0] _RAND_125;
  reg  _T_126; // @[Reg.scala 15:16]
  reg [31:0] _RAND_126;
  reg  _T_127; // @[Reg.scala 15:16]
  reg [31:0] _RAND_127;
  reg  _T_128; // @[Reg.scala 15:16]
  reg [31:0] _RAND_128;
  reg  _T_129; // @[Reg.scala 15:16]
  reg [31:0] _RAND_129;
  reg  _T_130; // @[Reg.scala 15:16]
  reg [31:0] _RAND_130;
  reg  _T_131; // @[Reg.scala 15:16]
  reg [31:0] _RAND_131;
  reg  _T_132; // @[Reg.scala 15:16]
  reg [31:0] _RAND_132;
  reg  _T_133; // @[Reg.scala 15:16]
  reg [31:0] _RAND_133;
  reg  _T_134; // @[Reg.scala 15:16]
  reg [31:0] _RAND_134;
  reg  _T_135; // @[Reg.scala 15:16]
  reg [31:0] _RAND_135;
  reg  _T_136; // @[Reg.scala 15:16]
  reg [31:0] _RAND_136;
  reg  _T_137; // @[Reg.scala 15:16]
  reg [31:0] _RAND_137;
  reg  _T_138; // @[Reg.scala 15:16]
  reg [31:0] _RAND_138;
  reg  _T_139; // @[Reg.scala 15:16]
  reg [31:0] _RAND_139;
  reg  _T_140; // @[Reg.scala 15:16]
  reg [31:0] _RAND_140;
  reg  _T_141; // @[Reg.scala 15:16]
  reg [31:0] _RAND_141;
  reg  _T_142; // @[Reg.scala 15:16]
  reg [31:0] _RAND_142;
  reg  _T_143; // @[Reg.scala 15:16]
  reg [31:0] _RAND_143;
  reg  _T_144; // @[Reg.scala 15:16]
  reg [31:0] _RAND_144;
  reg  _T_145; // @[Reg.scala 15:16]
  reg [31:0] _RAND_145;
  reg  _T_146; // @[Reg.scala 15:16]
  reg [31:0] _RAND_146;
  reg  _T_147; // @[Reg.scala 15:16]
  reg [31:0] _RAND_147;
  reg  _T_148; // @[Reg.scala 15:16]
  reg [31:0] _RAND_148;
  reg  _T_149; // @[Reg.scala 15:16]
  reg [31:0] _RAND_149;
  reg  _T_150; // @[Reg.scala 15:16]
  reg [31:0] _RAND_150;
  reg  _T_151; // @[Reg.scala 15:16]
  reg [31:0] _RAND_151;
  reg  _T_152; // @[Reg.scala 15:16]
  reg [31:0] _RAND_152;
  reg  _T_153; // @[Reg.scala 15:16]
  reg [31:0] _RAND_153;
  reg  _T_154; // @[Reg.scala 15:16]
  reg [31:0] _RAND_154;
  reg  _T_155; // @[Reg.scala 15:16]
  reg [31:0] _RAND_155;
  reg  _T_156; // @[Reg.scala 15:16]
  reg [31:0] _RAND_156;
  reg  _T_157; // @[Reg.scala 15:16]
  reg [31:0] _RAND_157;
  reg  _T_158; // @[Reg.scala 15:16]
  reg [31:0] _RAND_158;
  reg  _T_159; // @[Reg.scala 15:16]
  reg [31:0] _RAND_159;
  reg  _T_160; // @[Reg.scala 15:16]
  reg [31:0] _RAND_160;
  reg  _T_161; // @[Reg.scala 15:16]
  reg [31:0] _RAND_161;
  reg  _T_162; // @[Reg.scala 15:16]
  reg [31:0] _RAND_162;
  reg  _T_163; // @[Reg.scala 15:16]
  reg [31:0] _RAND_163;
  reg  _T_164; // @[Reg.scala 15:16]
  reg [31:0] _RAND_164;
  assign io_to_pes_0_sig_stat2trans = _T_14; // @[pe.scala 139:41]
  assign io_to_pes_0_out_ready = io_to_pes_1_in_ready; // @[pe.scala 143:38]
  assign io_to_pes_1_in_valid = io_to_pes_0_out_valid; // @[pe.scala 122:23]
  assign io_to_pes_1_in_bits = io_to_pes_0_out_bits; // @[pe.scala 122:23]
  assign io_to_pes_1_sig_stat2trans = _T_29; // @[pe.scala 139:41]
  assign io_to_pes_1_out_ready = io_to_pes_2_in_ready; // @[pe.scala 143:38]
  assign io_to_pes_2_in_valid = io_to_pes_1_out_valid; // @[pe.scala 122:23]
  assign io_to_pes_2_in_bits = io_to_pes_1_out_bits; // @[pe.scala 122:23]
  assign io_to_pes_2_sig_stat2trans = _T_44; // @[pe.scala 139:41]
  assign io_to_pes_2_out_ready = io_to_pes_3_in_ready; // @[pe.scala 143:38]
  assign io_to_pes_3_in_valid = io_to_pes_2_out_valid; // @[pe.scala 122:23]
  assign io_to_pes_3_in_bits = io_to_pes_2_out_bits; // @[pe.scala 122:23]
  assign io_to_pes_3_sig_stat2trans = _T_59; // @[pe.scala 139:41]
  assign io_to_pes_3_out_ready = io_to_pes_4_in_ready; // @[pe.scala 143:38]
  assign io_to_pes_4_in_valid = io_to_pes_3_out_valid; // @[pe.scala 122:23]
  assign io_to_pes_4_in_bits = io_to_pes_3_out_bits; // @[pe.scala 122:23]
  assign io_to_pes_4_sig_stat2trans = _T_74; // @[pe.scala 139:41]
  assign io_to_pes_4_out_ready = io_to_pes_5_in_ready; // @[pe.scala 143:38]
  assign io_to_pes_5_in_valid = io_to_pes_4_out_valid; // @[pe.scala 122:23]
  assign io_to_pes_5_in_bits = io_to_pes_4_out_bits; // @[pe.scala 122:23]
  assign io_to_pes_5_sig_stat2trans = _T_89; // @[pe.scala 139:41]
  assign io_to_pes_5_out_ready = io_to_pes_6_in_ready; // @[pe.scala 143:38]
  assign io_to_pes_6_in_valid = io_to_pes_5_out_valid; // @[pe.scala 122:23]
  assign io_to_pes_6_in_bits = io_to_pes_5_out_bits; // @[pe.scala 122:23]
  assign io_to_pes_6_sig_stat2trans = _T_104; // @[pe.scala 139:41]
  assign io_to_pes_6_out_ready = io_to_pes_7_in_ready; // @[pe.scala 143:38]
  assign io_to_pes_7_in_valid = io_to_pes_6_out_valid; // @[pe.scala 122:23]
  assign io_to_pes_7_in_bits = io_to_pes_6_out_bits; // @[pe.scala 122:23]
  assign io_to_pes_7_sig_stat2trans = _T_119; // @[pe.scala 139:41]
  assign io_to_pes_7_out_ready = io_to_pes_8_in_ready; // @[pe.scala 143:38]
  assign io_to_pes_8_in_valid = io_to_pes_7_out_valid; // @[pe.scala 122:23]
  assign io_to_pes_8_in_bits = io_to_pes_7_out_bits; // @[pe.scala 122:23]
  assign io_to_pes_8_sig_stat2trans = _T_134; // @[pe.scala 139:41]
  assign io_to_pes_8_out_ready = io_to_pes_9_in_ready; // @[pe.scala 143:38]
  assign io_to_pes_9_in_valid = io_to_pes_8_out_valid; // @[pe.scala 122:23]
  assign io_to_pes_9_in_bits = io_to_pes_8_out_bits; // @[pe.scala 122:23]
  assign io_to_pes_9_sig_stat2trans = _T_149; // @[pe.scala 139:41]
  assign io_to_pes_9_out_ready = io_to_pes_10_in_ready; // @[pe.scala 143:38]
  assign io_to_pes_10_in_valid = io_to_pes_9_out_valid; // @[pe.scala 122:23]
  assign io_to_pes_10_in_bits = io_to_pes_9_out_bits; // @[pe.scala 122:23]
  assign io_to_pes_10_sig_stat2trans = _T_164; // @[pe.scala 139:41]
  assign io_to_mem_valid = io_to_pes_10_out_valid; // @[pe.scala 129:17]
  assign io_to_mem_bits = io_to_pes_10_out_bits; // @[pe.scala 129:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_4 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_5 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_6 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_7 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_8 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_9 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_10 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_11 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_12 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_13 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_14 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_15 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_16 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_17 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_18 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_19 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_20 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_21 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_22 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_23 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_24 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_25 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_26 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_27 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_28 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_29 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_30 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_31 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_32 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_33 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_34 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_35 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_36 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_37 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_38 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_39 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_40 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_41 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_42 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_43 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_44 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_45 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_46 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_47 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_48 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_49 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_50 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_51 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _T_52 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _T_53 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T_54 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T_55 = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _T_56 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _T_57 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T_58 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T_59 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _T_60 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _T_61 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T_62 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T_63 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _T_64 = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _T_65 = _RAND_65[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _T_66 = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _T_67 = _RAND_67[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _T_68 = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  _T_69 = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _T_70 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _T_71 = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  _T_72 = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  _T_73 = _RAND_73[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _T_74 = _RAND_74[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _T_75 = _RAND_75[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  _T_76 = _RAND_76[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  _T_77 = _RAND_77[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  _T_78 = _RAND_78[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  _T_79 = _RAND_79[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  _T_80 = _RAND_80[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  _T_81 = _RAND_81[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _T_82 = _RAND_82[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _T_83 = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  _T_84 = _RAND_84[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  _T_85 = _RAND_85[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _T_86 = _RAND_86[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  _T_87 = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  _T_88 = _RAND_88[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  _T_89 = _RAND_89[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  _T_90 = _RAND_90[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  _T_91 = _RAND_91[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  _T_92 = _RAND_92[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  _T_93 = _RAND_93[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _T_94 = _RAND_94[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  _T_95 = _RAND_95[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  _T_96 = _RAND_96[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  _T_97 = _RAND_97[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  _T_98 = _RAND_98[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  _T_99 = _RAND_99[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  _T_100 = _RAND_100[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  _T_101 = _RAND_101[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  _T_102 = _RAND_102[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  _T_103 = _RAND_103[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  _T_104 = _RAND_104[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  _T_105 = _RAND_105[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  _T_106 = _RAND_106[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  _T_107 = _RAND_107[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  _T_108 = _RAND_108[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  _T_109 = _RAND_109[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  _T_110 = _RAND_110[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  _T_111 = _RAND_111[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  _T_112 = _RAND_112[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  _T_113 = _RAND_113[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  _T_114 = _RAND_114[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  _T_115 = _RAND_115[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  _T_116 = _RAND_116[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  _T_117 = _RAND_117[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  _T_118 = _RAND_118[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  _T_119 = _RAND_119[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  _T_120 = _RAND_120[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  _T_121 = _RAND_121[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  _T_122 = _RAND_122[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  _T_123 = _RAND_123[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  _T_124 = _RAND_124[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  _T_125 = _RAND_125[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  _T_126 = _RAND_126[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  _T_127 = _RAND_127[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  _T_128 = _RAND_128[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  _T_129 = _RAND_129[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  _T_130 = _RAND_130[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  _T_131 = _RAND_131[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  _T_132 = _RAND_132[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  _T_133 = _RAND_133[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  _T_134 = _RAND_134[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  _T_135 = _RAND_135[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  _T_136 = _RAND_136[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  _T_137 = _RAND_137[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  _T_138 = _RAND_138[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  _T_139 = _RAND_139[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  _T_140 = _RAND_140[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  _T_141 = _RAND_141[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  _T_142 = _RAND_142[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  _T_143 = _RAND_143[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  _T_144 = _RAND_144[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  _T_145 = _RAND_145[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  _T_146 = _RAND_146[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  _T_147 = _RAND_147[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  _T_148 = _RAND_148[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  _T_149 = _RAND_149[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  _T_150 = _RAND_150[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  _T_151 = _RAND_151[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  _T_152 = _RAND_152[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  _T_153 = _RAND_153[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  _T_154 = _RAND_154[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  _T_155 = _RAND_155[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  _T_156 = _RAND_156[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  _T_157 = _RAND_157[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  _T_158 = _RAND_158[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  _T_159 = _RAND_159[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  _T_160 = _RAND_160[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  _T_161 = _RAND_161[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  _T_162 = _RAND_162[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  _T_163 = _RAND_163[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  _T_164 = _RAND_164[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T <= io_sig_stat2trans;
    _T_1 <= _T;
    _T_2 <= _T_1;
    _T_3 <= _T_2;
    _T_4 <= _T_3;
    _T_5 <= _T_4;
    _T_6 <= _T_5;
    _T_7 <= _T_6;
    _T_8 <= _T_7;
    _T_9 <= _T_8;
    _T_10 <= _T_9;
    _T_11 <= _T_10;
    _T_12 <= _T_11;
    _T_13 <= _T_12;
    _T_14 <= _T_13;
    _T_15 <= io_sig_stat2trans;
    _T_16 <= _T_15;
    _T_17 <= _T_16;
    _T_18 <= _T_17;
    _T_19 <= _T_18;
    _T_20 <= _T_19;
    _T_21 <= _T_20;
    _T_22 <= _T_21;
    _T_23 <= _T_22;
    _T_24 <= _T_23;
    _T_25 <= _T_24;
    _T_26 <= _T_25;
    _T_27 <= _T_26;
    _T_28 <= _T_27;
    _T_29 <= _T_28;
    _T_30 <= io_sig_stat2trans;
    _T_31 <= _T_30;
    _T_32 <= _T_31;
    _T_33 <= _T_32;
    _T_34 <= _T_33;
    _T_35 <= _T_34;
    _T_36 <= _T_35;
    _T_37 <= _T_36;
    _T_38 <= _T_37;
    _T_39 <= _T_38;
    _T_40 <= _T_39;
    _T_41 <= _T_40;
    _T_42 <= _T_41;
    _T_43 <= _T_42;
    _T_44 <= _T_43;
    _T_45 <= io_sig_stat2trans;
    _T_46 <= _T_45;
    _T_47 <= _T_46;
    _T_48 <= _T_47;
    _T_49 <= _T_48;
    _T_50 <= _T_49;
    _T_51 <= _T_50;
    _T_52 <= _T_51;
    _T_53 <= _T_52;
    _T_54 <= _T_53;
    _T_55 <= _T_54;
    _T_56 <= _T_55;
    _T_57 <= _T_56;
    _T_58 <= _T_57;
    _T_59 <= _T_58;
    _T_60 <= io_sig_stat2trans;
    _T_61 <= _T_60;
    _T_62 <= _T_61;
    _T_63 <= _T_62;
    _T_64 <= _T_63;
    _T_65 <= _T_64;
    _T_66 <= _T_65;
    _T_67 <= _T_66;
    _T_68 <= _T_67;
    _T_69 <= _T_68;
    _T_70 <= _T_69;
    _T_71 <= _T_70;
    _T_72 <= _T_71;
    _T_73 <= _T_72;
    _T_74 <= _T_73;
    _T_75 <= io_sig_stat2trans;
    _T_76 <= _T_75;
    _T_77 <= _T_76;
    _T_78 <= _T_77;
    _T_79 <= _T_78;
    _T_80 <= _T_79;
    _T_81 <= _T_80;
    _T_82 <= _T_81;
    _T_83 <= _T_82;
    _T_84 <= _T_83;
    _T_85 <= _T_84;
    _T_86 <= _T_85;
    _T_87 <= _T_86;
    _T_88 <= _T_87;
    _T_89 <= _T_88;
    _T_90 <= io_sig_stat2trans;
    _T_91 <= _T_90;
    _T_92 <= _T_91;
    _T_93 <= _T_92;
    _T_94 <= _T_93;
    _T_95 <= _T_94;
    _T_96 <= _T_95;
    _T_97 <= _T_96;
    _T_98 <= _T_97;
    _T_99 <= _T_98;
    _T_100 <= _T_99;
    _T_101 <= _T_100;
    _T_102 <= _T_101;
    _T_103 <= _T_102;
    _T_104 <= _T_103;
    _T_105 <= io_sig_stat2trans;
    _T_106 <= _T_105;
    _T_107 <= _T_106;
    _T_108 <= _T_107;
    _T_109 <= _T_108;
    _T_110 <= _T_109;
    _T_111 <= _T_110;
    _T_112 <= _T_111;
    _T_113 <= _T_112;
    _T_114 <= _T_113;
    _T_115 <= _T_114;
    _T_116 <= _T_115;
    _T_117 <= _T_116;
    _T_118 <= _T_117;
    _T_119 <= _T_118;
    _T_120 <= io_sig_stat2trans;
    _T_121 <= _T_120;
    _T_122 <= _T_121;
    _T_123 <= _T_122;
    _T_124 <= _T_123;
    _T_125 <= _T_124;
    _T_126 <= _T_125;
    _T_127 <= _T_126;
    _T_128 <= _T_127;
    _T_129 <= _T_128;
    _T_130 <= _T_129;
    _T_131 <= _T_130;
    _T_132 <= _T_131;
    _T_133 <= _T_132;
    _T_134 <= _T_133;
    _T_135 <= io_sig_stat2trans;
    _T_136 <= _T_135;
    _T_137 <= _T_136;
    _T_138 <= _T_137;
    _T_139 <= _T_138;
    _T_140 <= _T_139;
    _T_141 <= _T_140;
    _T_142 <= _T_141;
    _T_143 <= _T_142;
    _T_144 <= _T_143;
    _T_145 <= _T_144;
    _T_146 <= _T_145;
    _T_147 <= _T_146;
    _T_148 <= _T_147;
    _T_149 <= _T_148;
    _T_150 <= io_sig_stat2trans;
    _T_151 <= _T_150;
    _T_152 <= _T_151;
    _T_153 <= _T_152;
    _T_154 <= _T_153;
    _T_155 <= _T_154;
    _T_156 <= _T_155;
    _T_157 <= _T_156;
    _T_158 <= _T_157;
    _T_159 <= _T_158;
    _T_160 <= _T_159;
    _T_161 <= _T_160;
    _T_162 <= _T_161;
    _T_163 <= _T_162;
    _T_164 <= _T_163;
  end
endmodule
module MultiDimMem(
  input         clock,
  input         reset,
  input         io_rd_addr_valid,
  input  [1:0]  io_rd_addr_bits_0,
  input  [1:0]  io_rd_addr_bits_1,
  input  [1:0]  io_rd_addr_bits_2,
  output        io_rd_data_valid,
  output [31:0] io_rd_data_bits,
  input         io_wr_addr_valid,
  input  [1:0]  io_wr_addr_bits_0,
  input  [1:0]  io_wr_addr_bits_1,
  input  [1:0]  io_wr_addr_bits_2,
  input         io_wr_data_valid,
  input  [31:0] io_wr_data_bits
);
  reg [32:0] mem [0:3071]; // @[mem.scala 116:24]
  reg [63:0] _RAND_0;
  wire [32:0] mem_mem_output_data; // @[mem.scala 116:24]
  wire [11:0] mem_mem_output_addr; // @[mem.scala 116:24]
  reg [63:0] _RAND_1;
  wire [32:0] mem__T_61_data; // @[mem.scala 116:24]
  wire [11:0] mem__T_61_addr; // @[mem.scala 116:24]
  wire  mem__T_61_mask; // @[mem.scala 116:24]
  wire  mem__T_61_en; // @[mem.scala 116:24]
  reg  mem_mem_output_en_pipe_0;
  reg [31:0] _RAND_2;
  reg [11:0] mem_mem_output_addr_pipe_0;
  reg [31:0] _RAND_3;
  reg  rd_addr_reg_valid; // @[mem.scala 117:28]
  reg [31:0] _RAND_4;
  reg [15:0] rd_addr_reg_bits_2; // @[mem.scala 117:28]
  reg [31:0] _RAND_5;
  reg [15:0] rd_addr_reg_bits_1; // @[mem.scala 117:28]
  reg [31:0] _RAND_6;
  reg [15:0] rd_addr_reg_bits_0; // @[mem.scala 117:28]
  reg [31:0] _RAND_7;
  wire [15:0] _T_8 = rd_addr_reg_bits_0 + 16'h1; // @[mem.scala 128:102]
  wire  _T_9 = 2'h1 == io_rd_addr_bits_0; // @[Mux.scala 68:19]
  wire  _T_11 = 2'h0 == io_rd_addr_bits_0; // @[Mux.scala 68:19]
  wire [15:0] _T_13 = rd_addr_reg_bits_1 + 16'hc; // @[mem.scala 128:102]
  wire  _T_14 = 2'h1 == io_rd_addr_bits_1; // @[Mux.scala 68:19]
  wire  _T_16 = 2'h0 == io_rd_addr_bits_1; // @[Mux.scala 68:19]
  wire [15:0] _T_18 = rd_addr_reg_bits_2 + 16'hc0; // @[mem.scala 128:102]
  wire  _T_19 = 2'h1 == io_rd_addr_bits_2; // @[Mux.scala 68:19]
  wire  _T_21 = 2'h0 == io_rd_addr_bits_2; // @[Mux.scala 68:19]
  wire [15:0] _T_23 = rd_addr_reg_bits_0 + rd_addr_reg_bits_1; // @[mem.scala 132:46]
  wire [15:0] mem_rd_addr = _T_23 + rd_addr_reg_bits_2; // @[mem.scala 132:46]
  reg  mem_req_valid; // @[mem.scala 139:30]
  reg [31:0] _RAND_8;
  reg  wr_addr_reg_valid; // @[mem.scala 142:28]
  reg [31:0] _RAND_9;
  reg [15:0] wr_addr_reg_bits_2; // @[mem.scala 142:28]
  reg [31:0] _RAND_10;
  reg [15:0] wr_addr_reg_bits_1; // @[mem.scala 142:28]
  reg [31:0] _RAND_11;
  reg [15:0] wr_addr_reg_bits_0; // @[mem.scala 142:28]
  reg [31:0] _RAND_12;
  wire [15:0] _T_40 = wr_addr_reg_bits_0 + 16'h1; // @[mem.scala 154:102]
  wire  _T_41 = 2'h1 == io_wr_addr_bits_0; // @[Mux.scala 68:19]
  wire  _T_43 = 2'h0 == io_wr_addr_bits_0; // @[Mux.scala 68:19]
  wire [15:0] _T_45 = wr_addr_reg_bits_1 + 16'hc; // @[mem.scala 154:102]
  wire  _T_46 = 2'h1 == io_wr_addr_bits_1; // @[Mux.scala 68:19]
  wire  _T_48 = 2'h0 == io_wr_addr_bits_1; // @[Mux.scala 68:19]
  wire [15:0] _T_50 = wr_addr_reg_bits_2 + 16'hc0; // @[mem.scala 154:102]
  wire  _T_51 = 2'h1 == io_wr_addr_bits_2; // @[Mux.scala 68:19]
  wire  _T_53 = 2'h0 == io_wr_addr_bits_2; // @[Mux.scala 68:19]
  reg  wr_data_reg_valid; // @[mem.scala 161:28]
  reg [31:0] _RAND_13;
  reg [31:0] wr_data_reg_bits; // @[mem.scala 161:28]
  reg [31:0] _RAND_14;
  wire [15:0] _T_56 = wr_addr_reg_bits_0 + wr_addr_reg_bits_1; // @[mem.scala 162:46]
  wire [15:0] mem_wr_addr = _T_56 + wr_addr_reg_bits_2; // @[mem.scala 162:46]
  wire [32:0] _GEN_9 = {wr_data_reg_valid, 32'h0}; // @[mem.scala 165:47]
  wire [63:0] _T_58 = {{31'd0}, _GEN_9}; // @[mem.scala 165:47]
  wire [63:0] _GEN_10 = {{32'd0}, wr_data_reg_bits}; // @[mem.scala 165:61]
  wire [63:0] _T_59 = _T_58 | _GEN_10; // @[mem.scala 165:61]
  wire  _T_63 = ~reset; // @[mem.scala 167:9]
  assign mem_mem_output_addr = mem_mem_output_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_mem_output_data = mem[mem_mem_output_addr]; // @[mem.scala 116:24]
  `else
  assign mem_mem_output_data = mem_mem_output_addr >= 12'hc00 ? _RAND_1[32:0] : mem[mem_mem_output_addr]; // @[mem.scala 116:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem__T_61_data = _T_59[32:0];
  assign mem__T_61_addr = mem_wr_addr[11:0];
  assign mem__T_61_mask = 1'h1;
  assign mem__T_61_en = wr_addr_reg_valid;
  assign io_rd_data_valid = mem_req_valid & mem_mem_output_data[32]; // @[mem.scala 140:20]
  assign io_rd_data_bits = mem_req_valid ? mem_mem_output_data[31:0] : 32'h0; // @[mem.scala 141:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3072; initvar = initvar+1)
    mem[initvar] = _RAND_0[32:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {2{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  mem_mem_output_en_pipe_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  mem_mem_output_addr_pipe_0 = _RAND_3[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  rd_addr_reg_valid = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  rd_addr_reg_bits_2 = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  rd_addr_reg_bits_1 = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  rd_addr_reg_bits_0 = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  mem_req_valid = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  wr_addr_reg_valid = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  wr_addr_reg_bits_2 = _RAND_10[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  wr_addr_reg_bits_1 = _RAND_11[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  wr_addr_reg_bits_0 = _RAND_12[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  wr_data_reg_valid = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  wr_data_reg_bits = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(mem__T_61_en & mem__T_61_mask) begin
      mem[mem__T_61_addr] <= mem__T_61_data; // @[mem.scala 116:24]
    end
    mem_mem_output_en_pipe_0 <= rd_addr_reg_valid;
    if (rd_addr_reg_valid) begin
      mem_mem_output_addr_pipe_0 <= mem_rd_addr[11:0];
    end
    if (reset) begin
      rd_addr_reg_valid <= 1'h0;
    end else begin
      rd_addr_reg_valid <= io_rd_addr_valid;
    end
    if (reset) begin
      rd_addr_reg_bits_2 <= 16'h0;
    end else if (_T_21) begin
      rd_addr_reg_bits_2 <= 16'h0;
    end else if (_T_19) begin
      rd_addr_reg_bits_2 <= _T_18;
    end
    if (reset) begin
      rd_addr_reg_bits_1 <= 16'h0;
    end else if (_T_16) begin
      rd_addr_reg_bits_1 <= 16'h0;
    end else if (_T_14) begin
      rd_addr_reg_bits_1 <= _T_13;
    end
    if (reset) begin
      rd_addr_reg_bits_0 <= 16'h0;
    end else if (_T_11) begin
      rd_addr_reg_bits_0 <= 16'h0;
    end else if (_T_9) begin
      rd_addr_reg_bits_0 <= _T_8;
    end
    if (reset) begin
      mem_req_valid <= 1'h0;
    end else begin
      mem_req_valid <= rd_addr_reg_valid;
    end
    if (reset) begin
      wr_addr_reg_valid <= 1'h0;
    end else begin
      wr_addr_reg_valid <= io_wr_addr_valid;
    end
    if (reset) begin
      wr_addr_reg_bits_2 <= 16'h0;
    end else if (_T_53) begin
      wr_addr_reg_bits_2 <= 16'h0;
    end else if (_T_51) begin
      wr_addr_reg_bits_2 <= _T_50;
    end
    if (reset) begin
      wr_addr_reg_bits_1 <= 16'h0;
    end else if (_T_48) begin
      wr_addr_reg_bits_1 <= 16'h0;
    end else if (_T_46) begin
      wr_addr_reg_bits_1 <= _T_45;
    end
    if (reset) begin
      wr_addr_reg_bits_0 <= 16'h0;
    end else if (_T_43) begin
      wr_addr_reg_bits_0 <= 16'h0;
    end else if (_T_41) begin
      wr_addr_reg_bits_0 <= _T_40;
    end
    if (reset) begin
      wr_data_reg_valid <= 1'h0;
    end else begin
      wr_data_reg_valid <= io_wr_data_valid;
    end
    if (reset) begin
      wr_data_reg_bits <= 32'h0;
    end else begin
      wr_data_reg_bits <= io_wr_data_bits;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_63) begin
          $fwrite(32'h80000002,"wr_addr:%d %d, wr_data: %d, rd_addr:%d %d, rd_data: %d %d\n",mem_wr_addr,wr_addr_reg_valid,wr_data_reg_bits,mem_rd_addr,rd_addr_reg_valid,io_rd_data_valid,io_rd_data_bits); // @[mem.scala 167:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module MemController(
  input         clock,
  input         reset,
  input         io_rd_valid,
  input         io_wr_valid,
  output        io_rd_data_valid,
  output [31:0] io_rd_data_bits,
  input         io_wr_data_valid,
  input  [31:0] io_wr_data_bits
);
  wire  MultiDimMem_clock; // @[mem.scala 31:19]
  wire  MultiDimMem_reset; // @[mem.scala 31:19]
  wire  MultiDimMem_io_rd_addr_valid; // @[mem.scala 31:19]
  wire [1:0] MultiDimMem_io_rd_addr_bits_0; // @[mem.scala 31:19]
  wire [1:0] MultiDimMem_io_rd_addr_bits_1; // @[mem.scala 31:19]
  wire [1:0] MultiDimMem_io_rd_addr_bits_2; // @[mem.scala 31:19]
  wire  MultiDimMem_io_rd_data_valid; // @[mem.scala 31:19]
  wire [31:0] MultiDimMem_io_rd_data_bits; // @[mem.scala 31:19]
  wire  MultiDimMem_io_wr_addr_valid; // @[mem.scala 31:19]
  wire [1:0] MultiDimMem_io_wr_addr_bits_0; // @[mem.scala 31:19]
  wire [1:0] MultiDimMem_io_wr_addr_bits_1; // @[mem.scala 31:19]
  wire [1:0] MultiDimMem_io_wr_addr_bits_2; // @[mem.scala 31:19]
  wire  MultiDimMem_io_wr_data_valid; // @[mem.scala 31:19]
  wire [31:0] MultiDimMem_io_wr_data_bits; // @[mem.scala 31:19]
  wire  MultiDimTime_clock; // @[mem.scala 32:23]
  wire  MultiDimTime_reset; // @[mem.scala 32:23]
  wire  MultiDimTime_io_in; // @[mem.scala 32:23]
  wire [1:0] MultiDimTime_io_out_0; // @[mem.scala 32:23]
  wire [1:0] MultiDimTime_io_out_1; // @[mem.scala 32:23]
  wire [1:0] MultiDimTime_io_out_2; // @[mem.scala 32:23]
  wire [15:0] MultiDimTime_io_index_0; // @[mem.scala 32:23]
  wire [15:0] MultiDimTime_io_index_1; // @[mem.scala 32:23]
  wire [15:0] MultiDimTime_io_index_2; // @[mem.scala 32:23]
  wire  MultiDimTime_1_clock; // @[mem.scala 33:23]
  wire  MultiDimTime_1_reset; // @[mem.scala 33:23]
  wire  MultiDimTime_1_io_in; // @[mem.scala 33:23]
  wire [1:0] MultiDimTime_1_io_out_0; // @[mem.scala 33:23]
  wire [1:0] MultiDimTime_1_io_out_1; // @[mem.scala 33:23]
  wire [1:0] MultiDimTime_1_io_out_2; // @[mem.scala 33:23]
  wire [15:0] MultiDimTime_1_io_index_0; // @[mem.scala 33:23]
  wire [15:0] MultiDimTime_1_io_index_1; // @[mem.scala 33:23]
  wire [15:0] MultiDimTime_1_io_index_2; // @[mem.scala 33:23]
  MultiDimMem MultiDimMem ( // @[mem.scala 31:19]
    .clock(MultiDimMem_clock),
    .reset(MultiDimMem_reset),
    .io_rd_addr_valid(MultiDimMem_io_rd_addr_valid),
    .io_rd_addr_bits_0(MultiDimMem_io_rd_addr_bits_0),
    .io_rd_addr_bits_1(MultiDimMem_io_rd_addr_bits_1),
    .io_rd_addr_bits_2(MultiDimMem_io_rd_addr_bits_2),
    .io_rd_data_valid(MultiDimMem_io_rd_data_valid),
    .io_rd_data_bits(MultiDimMem_io_rd_data_bits),
    .io_wr_addr_valid(MultiDimMem_io_wr_addr_valid),
    .io_wr_addr_bits_0(MultiDimMem_io_wr_addr_bits_0),
    .io_wr_addr_bits_1(MultiDimMem_io_wr_addr_bits_1),
    .io_wr_addr_bits_2(MultiDimMem_io_wr_addr_bits_2),
    .io_wr_data_valid(MultiDimMem_io_wr_data_valid),
    .io_wr_data_bits(MultiDimMem_io_wr_data_bits)
  );
  MultiDimTime MultiDimTime ( // @[mem.scala 32:23]
    .clock(MultiDimTime_clock),
    .reset(MultiDimTime_reset),
    .io_in(MultiDimTime_io_in),
    .io_out_0(MultiDimTime_io_out_0),
    .io_out_1(MultiDimTime_io_out_1),
    .io_out_2(MultiDimTime_io_out_2),
    .io_index_0(MultiDimTime_io_index_0),
    .io_index_1(MultiDimTime_io_index_1),
    .io_index_2(MultiDimTime_io_index_2)
  );
  MultiDimTime MultiDimTime_1 ( // @[mem.scala 33:23]
    .clock(MultiDimTime_1_clock),
    .reset(MultiDimTime_1_reset),
    .io_in(MultiDimTime_1_io_in),
    .io_out_0(MultiDimTime_1_io_out_0),
    .io_out_1(MultiDimTime_1_io_out_1),
    .io_out_2(MultiDimTime_1_io_out_2),
    .io_index_0(MultiDimTime_1_io_index_0),
    .io_index_1(MultiDimTime_1_io_index_1),
    .io_index_2(MultiDimTime_1_io_index_2)
  );
  assign io_rd_data_valid = MultiDimMem_io_rd_data_valid; // @[mem.scala 50:14]
  assign io_rd_data_bits = MultiDimMem_io_rd_data_bits; // @[mem.scala 50:14]
  assign MultiDimMem_clock = clock;
  assign MultiDimMem_reset = reset;
  assign MultiDimMem_io_rd_addr_valid = io_rd_valid; // @[mem.scala 47:21]
  assign MultiDimMem_io_rd_addr_bits_0 = MultiDimTime_1_io_out_0; // @[mem.scala 46:20]
  assign MultiDimMem_io_rd_addr_bits_1 = MultiDimTime_1_io_out_1; // @[mem.scala 46:20]
  assign MultiDimMem_io_rd_addr_bits_2 = MultiDimTime_1_io_out_2; // @[mem.scala 46:20]
  assign MultiDimMem_io_wr_addr_valid = io_wr_valid; // @[mem.scala 43:21]
  assign MultiDimMem_io_wr_addr_bits_0 = MultiDimTime_io_out_0; // @[mem.scala 42:20]
  assign MultiDimMem_io_wr_addr_bits_1 = MultiDimTime_io_out_1; // @[mem.scala 42:20]
  assign MultiDimMem_io_wr_addr_bits_2 = MultiDimTime_io_out_2; // @[mem.scala 42:20]
  assign MultiDimMem_io_wr_data_valid = io_wr_data_valid; // @[mem.scala 51:15]
  assign MultiDimMem_io_wr_data_bits = io_wr_data_bits; // @[mem.scala 51:15]
  assign MultiDimTime_clock = clock;
  assign MultiDimTime_reset = reset;
  assign MultiDimTime_io_in = io_wr_valid; // @[mem.scala 41:14]
  assign MultiDimTime_1_clock = clock;
  assign MultiDimTime_1_reset = reset;
  assign MultiDimTime_1_io_in = io_rd_valid; // @[mem.scala 45:14]
endmodule
module MultiDimMem_11(
  input          clock,
  input          reset,
  input          io_rd_addr_valid,
  input  [1:0]   io_rd_addr_bits_0,
  input  [1:0]   io_rd_addr_bits_1,
  input  [1:0]   io_rd_addr_bits_2,
  output         io_rd_data_valid,
  output [255:0] io_rd_data_bits,
  input          io_wr_addr_valid,
  input  [1:0]   io_wr_addr_bits_0,
  input  [1:0]   io_wr_addr_bits_1,
  input  [1:0]   io_wr_addr_bits_2,
  input          io_wr_data_valid,
  input  [255:0] io_wr_data_bits
);
  reg [256:0] mem [0:3071]; // @[mem.scala 116:24]
  reg [287:0] _RAND_0;
  wire [256:0] mem_mem_output_data; // @[mem.scala 116:24]
  wire [11:0] mem_mem_output_addr; // @[mem.scala 116:24]
  reg [287:0] _RAND_1;
  wire [256:0] mem__T_61_data; // @[mem.scala 116:24]
  wire [11:0] mem__T_61_addr; // @[mem.scala 116:24]
  wire  mem__T_61_mask; // @[mem.scala 116:24]
  wire  mem__T_61_en; // @[mem.scala 116:24]
  reg  mem_mem_output_en_pipe_0;
  reg [31:0] _RAND_2;
  reg [11:0] mem_mem_output_addr_pipe_0;
  reg [31:0] _RAND_3;
  reg  rd_addr_reg_valid; // @[mem.scala 117:28]
  reg [31:0] _RAND_4;
  reg [15:0] rd_addr_reg_bits_2; // @[mem.scala 117:28]
  reg [31:0] _RAND_5;
  reg [15:0] rd_addr_reg_bits_1; // @[mem.scala 117:28]
  reg [31:0] _RAND_6;
  reg [15:0] rd_addr_reg_bits_0; // @[mem.scala 117:28]
  reg [31:0] _RAND_7;
  wire [15:0] _T_8 = rd_addr_reg_bits_0 + 16'h1; // @[mem.scala 128:102]
  wire  _T_9 = 2'h1 == io_rd_addr_bits_0; // @[Mux.scala 68:19]
  wire  _T_11 = 2'h0 == io_rd_addr_bits_0; // @[Mux.scala 68:19]
  wire [15:0] _T_13 = rd_addr_reg_bits_1 + 16'hc; // @[mem.scala 128:102]
  wire  _T_14 = 2'h1 == io_rd_addr_bits_1; // @[Mux.scala 68:19]
  wire  _T_16 = 2'h0 == io_rd_addr_bits_1; // @[Mux.scala 68:19]
  wire [15:0] _T_18 = rd_addr_reg_bits_2 + 16'hc0; // @[mem.scala 128:102]
  wire  _T_19 = 2'h1 == io_rd_addr_bits_2; // @[Mux.scala 68:19]
  wire  _T_21 = 2'h0 == io_rd_addr_bits_2; // @[Mux.scala 68:19]
  wire [15:0] _T_23 = rd_addr_reg_bits_0 + rd_addr_reg_bits_1; // @[mem.scala 132:46]
  wire [15:0] mem_rd_addr = _T_23 + rd_addr_reg_bits_2; // @[mem.scala 132:46]
  reg  mem_req_valid; // @[mem.scala 139:30]
  reg [31:0] _RAND_8;
  reg  wr_addr_reg_valid; // @[mem.scala 142:28]
  reg [31:0] _RAND_9;
  reg [15:0] wr_addr_reg_bits_2; // @[mem.scala 142:28]
  reg [31:0] _RAND_10;
  reg [15:0] wr_addr_reg_bits_1; // @[mem.scala 142:28]
  reg [31:0] _RAND_11;
  reg [15:0] wr_addr_reg_bits_0; // @[mem.scala 142:28]
  reg [31:0] _RAND_12;
  wire [15:0] _T_40 = wr_addr_reg_bits_0 + 16'h1; // @[mem.scala 154:102]
  wire  _T_41 = 2'h1 == io_wr_addr_bits_0; // @[Mux.scala 68:19]
  wire  _T_43 = 2'h0 == io_wr_addr_bits_0; // @[Mux.scala 68:19]
  wire [15:0] _T_45 = wr_addr_reg_bits_1 + 16'hc; // @[mem.scala 154:102]
  wire  _T_46 = 2'h1 == io_wr_addr_bits_1; // @[Mux.scala 68:19]
  wire  _T_48 = 2'h0 == io_wr_addr_bits_1; // @[Mux.scala 68:19]
  wire [15:0] _T_50 = wr_addr_reg_bits_2 + 16'hc0; // @[mem.scala 154:102]
  wire  _T_51 = 2'h1 == io_wr_addr_bits_2; // @[Mux.scala 68:19]
  wire  _T_53 = 2'h0 == io_wr_addr_bits_2; // @[Mux.scala 68:19]
  reg  wr_data_reg_valid; // @[mem.scala 161:28]
  reg [31:0] _RAND_13;
  reg [255:0] wr_data_reg_bits; // @[mem.scala 161:28]
  reg [255:0] _RAND_14;
  wire [15:0] _T_56 = wr_addr_reg_bits_0 + wr_addr_reg_bits_1; // @[mem.scala 162:46]
  wire [15:0] mem_wr_addr = _T_56 + wr_addr_reg_bits_2; // @[mem.scala 162:46]
  wire [256:0] _GEN_9 = {wr_data_reg_valid, 256'h0}; // @[mem.scala 165:47]
  wire [511:0] _T_58 = {{255'd0}, _GEN_9}; // @[mem.scala 165:47]
  wire [511:0] _GEN_10 = {{256'd0}, wr_data_reg_bits}; // @[mem.scala 165:61]
  wire [511:0] _T_59 = _T_58 | _GEN_10; // @[mem.scala 165:61]
  wire  _T_63 = ~reset; // @[mem.scala 167:9]
  assign mem_mem_output_addr = mem_mem_output_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_mem_output_data = mem[mem_mem_output_addr]; // @[mem.scala 116:24]
  `else
  assign mem_mem_output_data = mem_mem_output_addr >= 12'hc00 ? _RAND_1[256:0] : mem[mem_mem_output_addr]; // @[mem.scala 116:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem__T_61_data = _T_59[256:0];
  assign mem__T_61_addr = mem_wr_addr[11:0];
  assign mem__T_61_mask = 1'h1;
  assign mem__T_61_en = wr_addr_reg_valid;
  assign io_rd_data_valid = mem_req_valid & mem_mem_output_data[256]; // @[mem.scala 140:20]
  assign io_rd_data_bits = mem_req_valid ? mem_mem_output_data[255:0] : 256'h0; // @[mem.scala 141:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {9{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 3072; initvar = initvar+1)
    mem[initvar] = _RAND_0[256:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {9{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  mem_mem_output_en_pipe_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  mem_mem_output_addr_pipe_0 = _RAND_3[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  rd_addr_reg_valid = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  rd_addr_reg_bits_2 = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  rd_addr_reg_bits_1 = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  rd_addr_reg_bits_0 = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  mem_req_valid = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  wr_addr_reg_valid = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  wr_addr_reg_bits_2 = _RAND_10[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  wr_addr_reg_bits_1 = _RAND_11[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  wr_addr_reg_bits_0 = _RAND_12[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  wr_data_reg_valid = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {8{`RANDOM}};
  wr_data_reg_bits = _RAND_14[255:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(mem__T_61_en & mem__T_61_mask) begin
      mem[mem__T_61_addr] <= mem__T_61_data; // @[mem.scala 116:24]
    end
    mem_mem_output_en_pipe_0 <= rd_addr_reg_valid;
    if (rd_addr_reg_valid) begin
      mem_mem_output_addr_pipe_0 <= mem_rd_addr[11:0];
    end
    if (reset) begin
      rd_addr_reg_valid <= 1'h0;
    end else begin
      rd_addr_reg_valid <= io_rd_addr_valid;
    end
    if (reset) begin
      rd_addr_reg_bits_2 <= 16'h0;
    end else if (_T_21) begin
      rd_addr_reg_bits_2 <= 16'h0;
    end else if (_T_19) begin
      rd_addr_reg_bits_2 <= _T_18;
    end
    if (reset) begin
      rd_addr_reg_bits_1 <= 16'h0;
    end else if (_T_16) begin
      rd_addr_reg_bits_1 <= 16'h0;
    end else if (_T_14) begin
      rd_addr_reg_bits_1 <= _T_13;
    end
    if (reset) begin
      rd_addr_reg_bits_0 <= 16'h0;
    end else if (_T_11) begin
      rd_addr_reg_bits_0 <= 16'h0;
    end else if (_T_9) begin
      rd_addr_reg_bits_0 <= _T_8;
    end
    if (reset) begin
      mem_req_valid <= 1'h0;
    end else begin
      mem_req_valid <= rd_addr_reg_valid;
    end
    if (reset) begin
      wr_addr_reg_valid <= 1'h0;
    end else begin
      wr_addr_reg_valid <= io_wr_addr_valid;
    end
    if (reset) begin
      wr_addr_reg_bits_2 <= 16'h0;
    end else if (_T_53) begin
      wr_addr_reg_bits_2 <= 16'h0;
    end else if (_T_51) begin
      wr_addr_reg_bits_2 <= _T_50;
    end
    if (reset) begin
      wr_addr_reg_bits_1 <= 16'h0;
    end else if (_T_48) begin
      wr_addr_reg_bits_1 <= 16'h0;
    end else if (_T_46) begin
      wr_addr_reg_bits_1 <= _T_45;
    end
    if (reset) begin
      wr_addr_reg_bits_0 <= 16'h0;
    end else if (_T_43) begin
      wr_addr_reg_bits_0 <= 16'h0;
    end else if (_T_41) begin
      wr_addr_reg_bits_0 <= _T_40;
    end
    if (reset) begin
      wr_data_reg_valid <= 1'h0;
    end else begin
      wr_data_reg_valid <= io_wr_data_valid;
    end
    if (reset) begin
      wr_data_reg_bits <= 256'h0;
    end else begin
      wr_data_reg_bits <= io_wr_data_bits;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_63) begin
          $fwrite(32'h80000002,"wr_addr:%d %d, wr_data: %d, rd_addr:%d %d, rd_data: %d %d\n",mem_wr_addr,wr_addr_reg_valid,wr_data_reg_bits,mem_rd_addr,rd_addr_reg_valid,io_rd_data_valid,io_rd_data_bits); // @[mem.scala 167:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module MemController_11(
  input          clock,
  input          reset,
  input          io_rd_valid,
  input          io_wr_valid,
  output         io_rd_data_valid,
  output [255:0] io_rd_data_bits,
  input          io_wr_data_valid,
  input  [255:0] io_wr_data_bits
);
  wire  MultiDimMem_clock; // @[mem.scala 31:19]
  wire  MultiDimMem_reset; // @[mem.scala 31:19]
  wire  MultiDimMem_io_rd_addr_valid; // @[mem.scala 31:19]
  wire [1:0] MultiDimMem_io_rd_addr_bits_0; // @[mem.scala 31:19]
  wire [1:0] MultiDimMem_io_rd_addr_bits_1; // @[mem.scala 31:19]
  wire [1:0] MultiDimMem_io_rd_addr_bits_2; // @[mem.scala 31:19]
  wire  MultiDimMem_io_rd_data_valid; // @[mem.scala 31:19]
  wire [255:0] MultiDimMem_io_rd_data_bits; // @[mem.scala 31:19]
  wire  MultiDimMem_io_wr_addr_valid; // @[mem.scala 31:19]
  wire [1:0] MultiDimMem_io_wr_addr_bits_0; // @[mem.scala 31:19]
  wire [1:0] MultiDimMem_io_wr_addr_bits_1; // @[mem.scala 31:19]
  wire [1:0] MultiDimMem_io_wr_addr_bits_2; // @[mem.scala 31:19]
  wire  MultiDimMem_io_wr_data_valid; // @[mem.scala 31:19]
  wire [255:0] MultiDimMem_io_wr_data_bits; // @[mem.scala 31:19]
  wire  MultiDimTime_clock; // @[mem.scala 32:23]
  wire  MultiDimTime_reset; // @[mem.scala 32:23]
  wire  MultiDimTime_io_in; // @[mem.scala 32:23]
  wire [1:0] MultiDimTime_io_out_0; // @[mem.scala 32:23]
  wire [1:0] MultiDimTime_io_out_1; // @[mem.scala 32:23]
  wire [1:0] MultiDimTime_io_out_2; // @[mem.scala 32:23]
  wire [15:0] MultiDimTime_io_index_0; // @[mem.scala 32:23]
  wire [15:0] MultiDimTime_io_index_1; // @[mem.scala 32:23]
  wire [15:0] MultiDimTime_io_index_2; // @[mem.scala 32:23]
  wire  MultiDimTime_1_clock; // @[mem.scala 33:23]
  wire  MultiDimTime_1_reset; // @[mem.scala 33:23]
  wire  MultiDimTime_1_io_in; // @[mem.scala 33:23]
  wire [1:0] MultiDimTime_1_io_out_0; // @[mem.scala 33:23]
  wire [1:0] MultiDimTime_1_io_out_1; // @[mem.scala 33:23]
  wire [1:0] MultiDimTime_1_io_out_2; // @[mem.scala 33:23]
  wire [15:0] MultiDimTime_1_io_index_0; // @[mem.scala 33:23]
  wire [15:0] MultiDimTime_1_io_index_1; // @[mem.scala 33:23]
  wire [15:0] MultiDimTime_1_io_index_2; // @[mem.scala 33:23]
  MultiDimMem_11 MultiDimMem ( // @[mem.scala 31:19]
    .clock(MultiDimMem_clock),
    .reset(MultiDimMem_reset),
    .io_rd_addr_valid(MultiDimMem_io_rd_addr_valid),
    .io_rd_addr_bits_0(MultiDimMem_io_rd_addr_bits_0),
    .io_rd_addr_bits_1(MultiDimMem_io_rd_addr_bits_1),
    .io_rd_addr_bits_2(MultiDimMem_io_rd_addr_bits_2),
    .io_rd_data_valid(MultiDimMem_io_rd_data_valid),
    .io_rd_data_bits(MultiDimMem_io_rd_data_bits),
    .io_wr_addr_valid(MultiDimMem_io_wr_addr_valid),
    .io_wr_addr_bits_0(MultiDimMem_io_wr_addr_bits_0),
    .io_wr_addr_bits_1(MultiDimMem_io_wr_addr_bits_1),
    .io_wr_addr_bits_2(MultiDimMem_io_wr_addr_bits_2),
    .io_wr_data_valid(MultiDimMem_io_wr_data_valid),
    .io_wr_data_bits(MultiDimMem_io_wr_data_bits)
  );
  MultiDimTime MultiDimTime ( // @[mem.scala 32:23]
    .clock(MultiDimTime_clock),
    .reset(MultiDimTime_reset),
    .io_in(MultiDimTime_io_in),
    .io_out_0(MultiDimTime_io_out_0),
    .io_out_1(MultiDimTime_io_out_1),
    .io_out_2(MultiDimTime_io_out_2),
    .io_index_0(MultiDimTime_io_index_0),
    .io_index_1(MultiDimTime_io_index_1),
    .io_index_2(MultiDimTime_io_index_2)
  );
  MultiDimTime MultiDimTime_1 ( // @[mem.scala 33:23]
    .clock(MultiDimTime_1_clock),
    .reset(MultiDimTime_1_reset),
    .io_in(MultiDimTime_1_io_in),
    .io_out_0(MultiDimTime_1_io_out_0),
    .io_out_1(MultiDimTime_1_io_out_1),
    .io_out_2(MultiDimTime_1_io_out_2),
    .io_index_0(MultiDimTime_1_io_index_0),
    .io_index_1(MultiDimTime_1_io_index_1),
    .io_index_2(MultiDimTime_1_io_index_2)
  );
  assign io_rd_data_valid = MultiDimMem_io_rd_data_valid; // @[mem.scala 50:14]
  assign io_rd_data_bits = MultiDimMem_io_rd_data_bits; // @[mem.scala 50:14]
  assign MultiDimMem_clock = clock;
  assign MultiDimMem_reset = reset;
  assign MultiDimMem_io_rd_addr_valid = io_rd_valid; // @[mem.scala 47:21]
  assign MultiDimMem_io_rd_addr_bits_0 = MultiDimTime_1_io_out_0; // @[mem.scala 46:20]
  assign MultiDimMem_io_rd_addr_bits_1 = MultiDimTime_1_io_out_1; // @[mem.scala 46:20]
  assign MultiDimMem_io_rd_addr_bits_2 = MultiDimTime_1_io_out_2; // @[mem.scala 46:20]
  assign MultiDimMem_io_wr_addr_valid = io_wr_valid; // @[mem.scala 43:21]
  assign MultiDimMem_io_wr_addr_bits_0 = MultiDimTime_io_out_0; // @[mem.scala 42:20]
  assign MultiDimMem_io_wr_addr_bits_1 = MultiDimTime_io_out_1; // @[mem.scala 42:20]
  assign MultiDimMem_io_wr_addr_bits_2 = MultiDimTime_io_out_2; // @[mem.scala 42:20]
  assign MultiDimMem_io_wr_data_valid = io_wr_data_valid; // @[mem.scala 51:15]
  assign MultiDimMem_io_wr_data_bits = io_wr_data_bits; // @[mem.scala 51:15]
  assign MultiDimTime_clock = clock;
  assign MultiDimTime_reset = reset;
  assign MultiDimTime_io_in = io_wr_valid; // @[mem.scala 41:14]
  assign MultiDimTime_1_clock = clock;
  assign MultiDimTime_1_reset = reset;
  assign MultiDimTime_1_io_in = io_rd_valid; // @[mem.scala 45:14]
endmodule
module MultiDimMem_26(
  input          clock,
  input          reset,
  input          io_rd_addr_valid,
  input  [1:0]   io_rd_addr_bits_0,
  input  [1:0]   io_rd_addr_bits_1,
  input  [1:0]   io_rd_addr_bits_2,
  output         io_rd_data_valid,
  output [255:0] io_rd_data_bits,
  input          io_wr_addr_valid,
  input  [1:0]   io_wr_addr_bits_0,
  input  [1:0]   io_wr_addr_bits_1,
  input  [1:0]   io_wr_addr_bits_2,
  input          io_wr_data_valid,
  input  [255:0] io_wr_data_bits
);
  reg [256:0] mem [0:2111]; // @[mem.scala 116:24]
  reg [287:0] _RAND_0;
  wire [256:0] mem_mem_output_data; // @[mem.scala 116:24]
  wire [11:0] mem_mem_output_addr; // @[mem.scala 116:24]
  reg [287:0] _RAND_1;
  wire [256:0] mem__T_61_data; // @[mem.scala 116:24]
  wire [11:0] mem__T_61_addr; // @[mem.scala 116:24]
  wire  mem__T_61_mask; // @[mem.scala 116:24]
  wire  mem__T_61_en; // @[mem.scala 116:24]
  reg  mem_mem_output_en_pipe_0;
  reg [31:0] _RAND_2;
  reg [11:0] mem_mem_output_addr_pipe_0;
  reg [31:0] _RAND_3;
  reg  rd_addr_reg_valid; // @[mem.scala 117:28]
  reg [31:0] _RAND_4;
  reg [15:0] rd_addr_reg_bits_2; // @[mem.scala 117:28]
  reg [31:0] _RAND_5;
  reg [15:0] rd_addr_reg_bits_1; // @[mem.scala 117:28]
  reg [31:0] _RAND_6;
  reg [15:0] rd_addr_reg_bits_0; // @[mem.scala 117:28]
  reg [31:0] _RAND_7;
  wire [15:0] _T_8 = rd_addr_reg_bits_0 + 16'h1; // @[mem.scala 128:102]
  wire  _T_9 = 2'h1 == io_rd_addr_bits_0; // @[Mux.scala 68:19]
  wire  _T_11 = 2'h0 == io_rd_addr_bits_0; // @[Mux.scala 68:19]
  wire [15:0] _T_13 = rd_addr_reg_bits_1 + 16'hc; // @[mem.scala 128:102]
  wire  _T_14 = 2'h1 == io_rd_addr_bits_1; // @[Mux.scala 68:19]
  wire  _T_16 = 2'h0 == io_rd_addr_bits_1; // @[Mux.scala 68:19]
  wire [15:0] _T_18 = rd_addr_reg_bits_2 + 16'h84; // @[mem.scala 128:102]
  wire  _T_19 = 2'h1 == io_rd_addr_bits_2; // @[Mux.scala 68:19]
  wire  _T_21 = 2'h0 == io_rd_addr_bits_2; // @[Mux.scala 68:19]
  wire [15:0] _T_23 = rd_addr_reg_bits_0 + rd_addr_reg_bits_1; // @[mem.scala 132:46]
  wire [15:0] mem_rd_addr = _T_23 + rd_addr_reg_bits_2; // @[mem.scala 132:46]
  reg  mem_req_valid; // @[mem.scala 139:30]
  reg [31:0] _RAND_8;
  reg  wr_addr_reg_valid; // @[mem.scala 142:28]
  reg [31:0] _RAND_9;
  reg [15:0] wr_addr_reg_bits_2; // @[mem.scala 142:28]
  reg [31:0] _RAND_10;
  reg [15:0] wr_addr_reg_bits_1; // @[mem.scala 142:28]
  reg [31:0] _RAND_11;
  reg [15:0] wr_addr_reg_bits_0; // @[mem.scala 142:28]
  reg [31:0] _RAND_12;
  wire [15:0] _T_40 = wr_addr_reg_bits_0 + 16'h1; // @[mem.scala 154:102]
  wire  _T_41 = 2'h1 == io_wr_addr_bits_0; // @[Mux.scala 68:19]
  wire  _T_43 = 2'h0 == io_wr_addr_bits_0; // @[Mux.scala 68:19]
  wire [15:0] _T_45 = wr_addr_reg_bits_1 + 16'hc; // @[mem.scala 154:102]
  wire  _T_46 = 2'h1 == io_wr_addr_bits_1; // @[Mux.scala 68:19]
  wire  _T_48 = 2'h0 == io_wr_addr_bits_1; // @[Mux.scala 68:19]
  wire [15:0] _T_50 = wr_addr_reg_bits_2 + 16'h84; // @[mem.scala 154:102]
  wire  _T_51 = 2'h1 == io_wr_addr_bits_2; // @[Mux.scala 68:19]
  wire  _T_53 = 2'h0 == io_wr_addr_bits_2; // @[Mux.scala 68:19]
  reg  wr_data_reg_valid; // @[mem.scala 161:28]
  reg [31:0] _RAND_13;
  reg [255:0] wr_data_reg_bits; // @[mem.scala 161:28]
  reg [255:0] _RAND_14;
  wire [15:0] _T_56 = wr_addr_reg_bits_0 + wr_addr_reg_bits_1; // @[mem.scala 162:46]
  wire [15:0] mem_wr_addr = _T_56 + wr_addr_reg_bits_2; // @[mem.scala 162:46]
  wire [256:0] _GEN_9 = {wr_data_reg_valid, 256'h0}; // @[mem.scala 165:47]
  wire [511:0] _T_58 = {{255'd0}, _GEN_9}; // @[mem.scala 165:47]
  wire [511:0] _GEN_10 = {{256'd0}, wr_data_reg_bits}; // @[mem.scala 165:61]
  wire [511:0] _T_59 = _T_58 | _GEN_10; // @[mem.scala 165:61]
  wire  _T_63 = ~reset; // @[mem.scala 167:9]
  assign mem_mem_output_addr = mem_mem_output_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign mem_mem_output_data = mem[mem_mem_output_addr]; // @[mem.scala 116:24]
  `else
  assign mem_mem_output_data = mem_mem_output_addr >= 12'h840 ? _RAND_1[256:0] : mem[mem_mem_output_addr]; // @[mem.scala 116:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign mem__T_61_data = _T_59[256:0];
  assign mem__T_61_addr = mem_wr_addr[11:0];
  assign mem__T_61_mask = 1'h1;
  assign mem__T_61_en = wr_addr_reg_valid;
  assign io_rd_data_valid = mem_req_valid & mem_mem_output_data[256]; // @[mem.scala 140:20]
  assign io_rd_data_bits = mem_req_valid ? mem_mem_output_data[255:0] : 256'h0; // @[mem.scala 141:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {9{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2112; initvar = initvar+1)
    mem[initvar] = _RAND_0[256:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {9{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  mem_mem_output_en_pipe_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  mem_mem_output_addr_pipe_0 = _RAND_3[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  rd_addr_reg_valid = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  rd_addr_reg_bits_2 = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  rd_addr_reg_bits_1 = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  rd_addr_reg_bits_0 = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  mem_req_valid = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  wr_addr_reg_valid = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  wr_addr_reg_bits_2 = _RAND_10[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  wr_addr_reg_bits_1 = _RAND_11[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  wr_addr_reg_bits_0 = _RAND_12[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  wr_data_reg_valid = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {8{`RANDOM}};
  wr_data_reg_bits = _RAND_14[255:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(mem__T_61_en & mem__T_61_mask) begin
      mem[mem__T_61_addr] <= mem__T_61_data; // @[mem.scala 116:24]
    end
    mem_mem_output_en_pipe_0 <= rd_addr_reg_valid;
    if (rd_addr_reg_valid) begin
      mem_mem_output_addr_pipe_0 <= mem_rd_addr[11:0];
    end
    if (reset) begin
      rd_addr_reg_valid <= 1'h0;
    end else begin
      rd_addr_reg_valid <= io_rd_addr_valid;
    end
    if (reset) begin
      rd_addr_reg_bits_2 <= 16'h0;
    end else if (_T_21) begin
      rd_addr_reg_bits_2 <= 16'h0;
    end else if (_T_19) begin
      rd_addr_reg_bits_2 <= _T_18;
    end
    if (reset) begin
      rd_addr_reg_bits_1 <= 16'h0;
    end else if (_T_16) begin
      rd_addr_reg_bits_1 <= 16'h0;
    end else if (_T_14) begin
      rd_addr_reg_bits_1 <= _T_13;
    end
    if (reset) begin
      rd_addr_reg_bits_0 <= 16'h0;
    end else if (_T_11) begin
      rd_addr_reg_bits_0 <= 16'h0;
    end else if (_T_9) begin
      rd_addr_reg_bits_0 <= _T_8;
    end
    if (reset) begin
      mem_req_valid <= 1'h0;
    end else begin
      mem_req_valid <= rd_addr_reg_valid;
    end
    if (reset) begin
      wr_addr_reg_valid <= 1'h0;
    end else begin
      wr_addr_reg_valid <= io_wr_addr_valid;
    end
    if (reset) begin
      wr_addr_reg_bits_2 <= 16'h0;
    end else if (_T_53) begin
      wr_addr_reg_bits_2 <= 16'h0;
    end else if (_T_51) begin
      wr_addr_reg_bits_2 <= _T_50;
    end
    if (reset) begin
      wr_addr_reg_bits_1 <= 16'h0;
    end else if (_T_48) begin
      wr_addr_reg_bits_1 <= 16'h0;
    end else if (_T_46) begin
      wr_addr_reg_bits_1 <= _T_45;
    end
    if (reset) begin
      wr_addr_reg_bits_0 <= 16'h0;
    end else if (_T_43) begin
      wr_addr_reg_bits_0 <= 16'h0;
    end else if (_T_41) begin
      wr_addr_reg_bits_0 <= _T_40;
    end
    if (reset) begin
      wr_data_reg_valid <= 1'h0;
    end else begin
      wr_data_reg_valid <= io_wr_data_valid;
    end
    if (reset) begin
      wr_data_reg_bits <= 256'h0;
    end else begin
      wr_data_reg_bits <= io_wr_data_bits;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_63) begin
          $fwrite(32'h80000002,"wr_addr:%d %d, wr_data: %d, rd_addr:%d %d, rd_data: %d %d\n",mem_wr_addr,wr_addr_reg_valid,wr_data_reg_bits,mem_rd_addr,rd_addr_reg_valid,io_rd_data_valid,io_rd_data_bits); // @[mem.scala 167:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module MultiDimTime_53(
  input        clock,
  input        reset,
  input        io_in,
  output [1:0] io_out_0,
  output [1:0] io_out_1,
  output [1:0] io_out_2
);
  reg [15:0] regs_0; // @[mem.scala 67:12]
  reg [31:0] _RAND_0;
  reg [15:0] regs_1; // @[mem.scala 67:12]
  reg [31:0] _RAND_1;
  reg [15:0] regs_2; // @[mem.scala 67:12]
  reg [31:0] _RAND_2;
  wire [15:0] _GEN_10 = {{15'd0}, io_in}; // @[mem.scala 69:42]
  wire [15:0] _T_1 = regs_0 + _GEN_10; // @[mem.scala 69:42]
  wire  back_0 = _T_1 == 16'hc; // @[mem.scala 69:48]
  wire [15:0] _T_3 = regs_1 + _GEN_10; // @[mem.scala 69:42]
  wire  next_1 = _T_3 == 16'hb; // @[mem.scala 69:48]
  wire [15:0] _T_5 = regs_2 + _GEN_10; // @[mem.scala 69:42]
  wire  next_2 = _T_5 == 16'h10; // @[mem.scala 69:48]
  wire  back_1 = back_0 & next_1; // @[mem.scala 71:32]
  wire  back_2 = back_1 & next_2; // @[mem.scala 71:32]
  wire  _GEN_1 = back_0 ? 1'h0 : io_in; // @[mem.scala 90:20]
  wire  _GEN_3 = back_1 ? 1'h0 : 1'h1; // @[mem.scala 79:22]
  wire  _GEN_7 = back_2 ? 1'h0 : 1'h1; // @[mem.scala 79:22]
  assign io_out_0 = {{1'd0}, _GEN_1}; // @[mem.scala 92:19 mem.scala 95:19]
  assign io_out_1 = back_0 ? {{1'd0}, _GEN_3} : 2'h2; // @[mem.scala 81:21 mem.scala 84:21 mem.scala 87:19]
  assign io_out_2 = back_1 ? {{1'd0}, _GEN_7} : 2'h2; // @[mem.scala 81:21 mem.scala 84:21 mem.scala 87:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 16'h0;
    end else if (back_0) begin
      regs_0 <= 16'h0;
    end else begin
      regs_0 <= _T_1;
    end
    if (reset) begin
      regs_1 <= 16'h0;
    end else if (back_0) begin
      if (back_1) begin
        regs_1 <= 16'h0;
      end else begin
        regs_1 <= _T_3;
      end
    end
    if (reset) begin
      regs_2 <= 16'h0;
    end else if (back_1) begin
      if (back_2) begin
        regs_2 <= 16'h0;
      end else begin
        regs_2 <= _T_5;
      end
    end
  end
endmodule
module MemController_26(
  input          clock,
  input          reset,
  input          io_rd_valid,
  input          io_wr_valid,
  output         io_rd_data_valid,
  output [255:0] io_rd_data_bits,
  input          io_wr_data_valid,
  input  [255:0] io_wr_data_bits
);
  wire  MultiDimMem_clock; // @[mem.scala 31:19]
  wire  MultiDimMem_reset; // @[mem.scala 31:19]
  wire  MultiDimMem_io_rd_addr_valid; // @[mem.scala 31:19]
  wire [1:0] MultiDimMem_io_rd_addr_bits_0; // @[mem.scala 31:19]
  wire [1:0] MultiDimMem_io_rd_addr_bits_1; // @[mem.scala 31:19]
  wire [1:0] MultiDimMem_io_rd_addr_bits_2; // @[mem.scala 31:19]
  wire  MultiDimMem_io_rd_data_valid; // @[mem.scala 31:19]
  wire [255:0] MultiDimMem_io_rd_data_bits; // @[mem.scala 31:19]
  wire  MultiDimMem_io_wr_addr_valid; // @[mem.scala 31:19]
  wire [1:0] MultiDimMem_io_wr_addr_bits_0; // @[mem.scala 31:19]
  wire [1:0] MultiDimMem_io_wr_addr_bits_1; // @[mem.scala 31:19]
  wire [1:0] MultiDimMem_io_wr_addr_bits_2; // @[mem.scala 31:19]
  wire  MultiDimMem_io_wr_data_valid; // @[mem.scala 31:19]
  wire [255:0] MultiDimMem_io_wr_data_bits; // @[mem.scala 31:19]
  wire  MultiDimTime_clock; // @[mem.scala 32:23]
  wire  MultiDimTime_reset; // @[mem.scala 32:23]
  wire  MultiDimTime_io_in; // @[mem.scala 32:23]
  wire [1:0] MultiDimTime_io_out_0; // @[mem.scala 32:23]
  wire [1:0] MultiDimTime_io_out_1; // @[mem.scala 32:23]
  wire [1:0] MultiDimTime_io_out_2; // @[mem.scala 32:23]
  wire  MultiDimTime_1_clock; // @[mem.scala 33:23]
  wire  MultiDimTime_1_reset; // @[mem.scala 33:23]
  wire  MultiDimTime_1_io_in; // @[mem.scala 33:23]
  wire [1:0] MultiDimTime_1_io_out_0; // @[mem.scala 33:23]
  wire [1:0] MultiDimTime_1_io_out_1; // @[mem.scala 33:23]
  wire [1:0] MultiDimTime_1_io_out_2; // @[mem.scala 33:23]
  MultiDimMem_26 MultiDimMem ( // @[mem.scala 31:19]
    .clock(MultiDimMem_clock),
    .reset(MultiDimMem_reset),
    .io_rd_addr_valid(MultiDimMem_io_rd_addr_valid),
    .io_rd_addr_bits_0(MultiDimMem_io_rd_addr_bits_0),
    .io_rd_addr_bits_1(MultiDimMem_io_rd_addr_bits_1),
    .io_rd_addr_bits_2(MultiDimMem_io_rd_addr_bits_2),
    .io_rd_data_valid(MultiDimMem_io_rd_data_valid),
    .io_rd_data_bits(MultiDimMem_io_rd_data_bits),
    .io_wr_addr_valid(MultiDimMem_io_wr_addr_valid),
    .io_wr_addr_bits_0(MultiDimMem_io_wr_addr_bits_0),
    .io_wr_addr_bits_1(MultiDimMem_io_wr_addr_bits_1),
    .io_wr_addr_bits_2(MultiDimMem_io_wr_addr_bits_2),
    .io_wr_data_valid(MultiDimMem_io_wr_data_valid),
    .io_wr_data_bits(MultiDimMem_io_wr_data_bits)
  );
  MultiDimTime_53 MultiDimTime ( // @[mem.scala 32:23]
    .clock(MultiDimTime_clock),
    .reset(MultiDimTime_reset),
    .io_in(MultiDimTime_io_in),
    .io_out_0(MultiDimTime_io_out_0),
    .io_out_1(MultiDimTime_io_out_1),
    .io_out_2(MultiDimTime_io_out_2)
  );
  MultiDimTime_53 MultiDimTime_1 ( // @[mem.scala 33:23]
    .clock(MultiDimTime_1_clock),
    .reset(MultiDimTime_1_reset),
    .io_in(MultiDimTime_1_io_in),
    .io_out_0(MultiDimTime_1_io_out_0),
    .io_out_1(MultiDimTime_1_io_out_1),
    .io_out_2(MultiDimTime_1_io_out_2)
  );
  assign io_rd_data_valid = MultiDimMem_io_rd_data_valid; // @[mem.scala 50:14]
  assign io_rd_data_bits = MultiDimMem_io_rd_data_bits; // @[mem.scala 50:14]
  assign MultiDimMem_clock = clock;
  assign MultiDimMem_reset = reset;
  assign MultiDimMem_io_rd_addr_valid = io_rd_valid; // @[mem.scala 47:21]
  assign MultiDimMem_io_rd_addr_bits_0 = MultiDimTime_1_io_out_0; // @[mem.scala 46:20]
  assign MultiDimMem_io_rd_addr_bits_1 = MultiDimTime_1_io_out_1; // @[mem.scala 46:20]
  assign MultiDimMem_io_rd_addr_bits_2 = MultiDimTime_1_io_out_2; // @[mem.scala 46:20]
  assign MultiDimMem_io_wr_addr_valid = io_wr_valid; // @[mem.scala 43:21]
  assign MultiDimMem_io_wr_addr_bits_0 = MultiDimTime_io_out_0; // @[mem.scala 42:20]
  assign MultiDimMem_io_wr_addr_bits_1 = MultiDimTime_io_out_1; // @[mem.scala 42:20]
  assign MultiDimMem_io_wr_addr_bits_2 = MultiDimTime_io_out_2; // @[mem.scala 42:20]
  assign MultiDimMem_io_wr_data_valid = io_wr_data_valid; // @[mem.scala 51:15]
  assign MultiDimMem_io_wr_data_bits = io_wr_data_bits; // @[mem.scala 51:15]
  assign MultiDimTime_clock = clock;
  assign MultiDimTime_reset = reset;
  assign MultiDimTime_io_in = io_wr_valid; // @[mem.scala 41:14]
  assign MultiDimTime_1_clock = clock;
  assign MultiDimTime_1_reset = reset;
  assign MultiDimTime_1_io_in = io_rd_valid; // @[mem.scala 45:14]
endmodule
module PEArray2D(
  input          clock,
  input          reset,
  output         io_data_2_out_0_valid,
  output [255:0] io_data_2_out_0_bits,
  output         io_data_2_out_1_valid,
  output [255:0] io_data_2_out_1_bits,
  output         io_data_2_out_2_valid,
  output [255:0] io_data_2_out_2_bits,
  output         io_data_2_out_3_valid,
  output [255:0] io_data_2_out_3_bits,
  output         io_data_2_out_4_valid,
  output [255:0] io_data_2_out_4_bits,
  output         io_data_2_out_5_valid,
  output [255:0] io_data_2_out_5_bits,
  output         io_data_2_out_6_valid,
  output [255:0] io_data_2_out_6_bits,
  output         io_data_2_out_7_valid,
  output [255:0] io_data_2_out_7_bits,
  output         io_data_2_out_8_valid,
  output [255:0] io_data_2_out_8_bits,
  output         io_data_2_out_9_valid,
  output [255:0] io_data_2_out_9_bits,
  output         io_data_2_out_10_valid,
  output [255:0] io_data_2_out_10_bits,
  output         io_data_2_out_11_valid,
  output [255:0] io_data_2_out_11_bits,
  output         io_data_2_out_12_valid,
  output [255:0] io_data_2_out_12_bits,
  output         io_data_2_out_13_valid,
  output [255:0] io_data_2_out_13_bits,
  output         io_data_2_out_14_valid,
  output [255:0] io_data_2_out_14_bits,
  input          io_data_1_in_0_valid,
  input          io_data_1_in_0_bits_valid,
  input  [255:0] io_data_1_in_0_bits_bits,
  input          io_data_1_in_1_valid,
  input          io_data_1_in_1_bits_valid,
  input  [255:0] io_data_1_in_1_bits_bits,
  input          io_data_1_in_2_valid,
  input          io_data_1_in_2_bits_valid,
  input  [255:0] io_data_1_in_2_bits_bits,
  input          io_data_1_in_3_valid,
  input          io_data_1_in_3_bits_valid,
  input  [255:0] io_data_1_in_3_bits_bits,
  input          io_data_1_in_4_valid,
  input          io_data_1_in_4_bits_valid,
  input  [255:0] io_data_1_in_4_bits_bits,
  input          io_data_1_in_5_valid,
  input          io_data_1_in_5_bits_valid,
  input  [255:0] io_data_1_in_5_bits_bits,
  input          io_data_1_in_6_valid,
  input          io_data_1_in_6_bits_valid,
  input  [255:0] io_data_1_in_6_bits_bits,
  input          io_data_1_in_7_valid,
  input          io_data_1_in_7_bits_valid,
  input  [255:0] io_data_1_in_7_bits_bits,
  input          io_data_1_in_8_valid,
  input          io_data_1_in_8_bits_valid,
  input  [255:0] io_data_1_in_8_bits_bits,
  input          io_data_1_in_9_valid,
  input          io_data_1_in_9_bits_valid,
  input  [255:0] io_data_1_in_9_bits_bits,
  input          io_data_1_in_10_valid,
  input          io_data_1_in_10_bits_valid,
  input  [255:0] io_data_1_in_10_bits_bits,
  input          io_data_1_in_11_valid,
  input          io_data_1_in_11_bits_valid,
  input  [255:0] io_data_1_in_11_bits_bits,
  input          io_data_1_in_12_valid,
  input          io_data_1_in_12_bits_valid,
  input  [255:0] io_data_1_in_12_bits_bits,
  input          io_data_1_in_13_valid,
  input          io_data_1_in_13_bits_valid,
  input  [255:0] io_data_1_in_13_bits_bits,
  input          io_data_1_in_14_valid,
  input          io_data_1_in_14_bits_valid,
  input  [255:0] io_data_1_in_14_bits_bits,
  input          io_data_0_in_0_valid,
  input          io_data_0_in_0_bits_valid,
  input  [31:0]  io_data_0_in_0_bits_bits,
  input          io_data_0_in_1_valid,
  input          io_data_0_in_1_bits_valid,
  input  [31:0]  io_data_0_in_1_bits_bits,
  input          io_data_0_in_2_valid,
  input          io_data_0_in_2_bits_valid,
  input  [31:0]  io_data_0_in_2_bits_bits,
  input          io_data_0_in_3_valid,
  input          io_data_0_in_3_bits_valid,
  input  [31:0]  io_data_0_in_3_bits_bits,
  input          io_data_0_in_4_valid,
  input          io_data_0_in_4_bits_valid,
  input  [31:0]  io_data_0_in_4_bits_bits,
  input          io_data_0_in_5_valid,
  input          io_data_0_in_5_bits_valid,
  input  [31:0]  io_data_0_in_5_bits_bits,
  input          io_data_0_in_6_valid,
  input          io_data_0_in_6_bits_valid,
  input  [31:0]  io_data_0_in_6_bits_bits,
  input          io_data_0_in_7_valid,
  input          io_data_0_in_7_bits_valid,
  input  [31:0]  io_data_0_in_7_bits_bits,
  input          io_data_0_in_8_valid,
  input          io_data_0_in_8_bits_valid,
  input  [31:0]  io_data_0_in_8_bits_bits,
  input          io_data_0_in_9_valid,
  input          io_data_0_in_9_bits_valid,
  input  [31:0]  io_data_0_in_9_bits_bits,
  input          io_data_0_in_10_valid,
  input          io_data_0_in_10_bits_valid,
  input  [31:0]  io_data_0_in_10_bits_bits,
  input          io_exec_valid,
  input          io_out_valid
);
  wire  MultiDimTime_clock; // @[pe.scala 162:25]
  wire  MultiDimTime_reset; // @[pe.scala 162:25]
  wire  MultiDimTime_io_in; // @[pe.scala 162:25]
  wire [1:0] MultiDimTime_io_out_0; // @[pe.scala 162:25]
  wire [1:0] MultiDimTime_io_out_1; // @[pe.scala 162:25]
  wire [1:0] MultiDimTime_io_out_2; // @[pe.scala 162:25]
  wire [15:0] MultiDimTime_io_index_0; // @[pe.scala 162:25]
  wire [15:0] MultiDimTime_io_index_1; // @[pe.scala 162:25]
  wire [15:0] MultiDimTime_io_index_2; // @[pe.scala 162:25]
  wire  PE_clock; // @[pe.scala 184:13]
  wire  PE_reset; // @[pe.scala 184:13]
  wire  PE_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_1_clock; // @[pe.scala 184:13]
  wire  PE_1_reset; // @[pe.scala 184:13]
  wire  PE_1_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_1_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_1_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_1_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_1_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_1_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_1_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_1_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_1_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_1_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_1_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_1_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_1_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_1_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_1_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_2_clock; // @[pe.scala 184:13]
  wire  PE_2_reset; // @[pe.scala 184:13]
  wire  PE_2_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_2_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_2_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_2_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_2_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_2_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_2_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_2_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_2_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_2_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_2_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_2_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_2_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_2_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_2_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_3_clock; // @[pe.scala 184:13]
  wire  PE_3_reset; // @[pe.scala 184:13]
  wire  PE_3_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_3_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_3_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_3_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_3_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_3_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_3_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_3_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_3_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_3_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_3_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_3_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_3_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_3_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_3_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_4_clock; // @[pe.scala 184:13]
  wire  PE_4_reset; // @[pe.scala 184:13]
  wire  PE_4_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_4_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_4_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_4_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_4_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_4_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_4_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_4_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_4_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_4_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_4_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_4_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_4_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_4_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_4_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_5_clock; // @[pe.scala 184:13]
  wire  PE_5_reset; // @[pe.scala 184:13]
  wire  PE_5_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_5_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_5_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_5_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_5_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_5_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_5_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_5_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_5_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_5_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_5_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_5_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_5_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_5_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_5_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_6_clock; // @[pe.scala 184:13]
  wire  PE_6_reset; // @[pe.scala 184:13]
  wire  PE_6_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_6_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_6_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_6_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_6_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_6_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_6_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_6_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_6_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_6_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_6_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_6_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_6_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_6_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_6_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_7_clock; // @[pe.scala 184:13]
  wire  PE_7_reset; // @[pe.scala 184:13]
  wire  PE_7_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_7_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_7_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_7_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_7_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_7_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_7_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_7_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_7_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_7_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_7_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_7_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_7_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_7_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_7_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_8_clock; // @[pe.scala 184:13]
  wire  PE_8_reset; // @[pe.scala 184:13]
  wire  PE_8_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_8_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_8_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_8_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_8_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_8_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_8_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_8_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_8_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_8_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_8_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_8_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_8_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_8_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_8_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_9_clock; // @[pe.scala 184:13]
  wire  PE_9_reset; // @[pe.scala 184:13]
  wire  PE_9_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_9_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_9_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_9_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_9_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_9_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_9_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_9_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_9_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_9_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_9_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_9_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_9_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_9_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_9_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_10_clock; // @[pe.scala 184:13]
  wire  PE_10_reset; // @[pe.scala 184:13]
  wire  PE_10_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_10_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_10_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_10_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_10_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_10_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_10_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_10_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_10_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_10_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_10_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_10_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_10_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_10_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_10_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_11_clock; // @[pe.scala 184:13]
  wire  PE_11_reset; // @[pe.scala 184:13]
  wire  PE_11_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_11_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_11_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_11_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_11_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_11_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_11_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_11_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_11_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_11_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_11_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_11_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_11_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_11_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_11_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_12_clock; // @[pe.scala 184:13]
  wire  PE_12_reset; // @[pe.scala 184:13]
  wire  PE_12_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_12_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_12_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_12_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_12_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_12_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_12_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_12_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_12_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_12_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_12_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_12_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_12_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_12_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_12_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_13_clock; // @[pe.scala 184:13]
  wire  PE_13_reset; // @[pe.scala 184:13]
  wire  PE_13_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_13_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_13_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_13_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_13_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_13_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_13_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_13_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_13_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_13_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_13_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_13_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_13_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_13_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_13_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_14_clock; // @[pe.scala 184:13]
  wire  PE_14_reset; // @[pe.scala 184:13]
  wire  PE_14_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_14_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_14_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_14_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_14_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_14_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_14_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_14_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_14_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_14_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_14_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_14_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_14_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_14_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_14_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_15_clock; // @[pe.scala 184:13]
  wire  PE_15_reset; // @[pe.scala 184:13]
  wire  PE_15_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_15_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_15_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_15_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_15_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_15_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_15_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_15_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_15_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_15_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_15_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_15_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_15_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_15_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_15_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_16_clock; // @[pe.scala 184:13]
  wire  PE_16_reset; // @[pe.scala 184:13]
  wire  PE_16_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_16_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_16_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_16_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_16_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_16_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_16_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_16_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_16_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_16_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_16_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_16_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_16_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_16_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_16_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_17_clock; // @[pe.scala 184:13]
  wire  PE_17_reset; // @[pe.scala 184:13]
  wire  PE_17_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_17_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_17_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_17_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_17_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_17_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_17_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_17_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_17_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_17_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_17_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_17_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_17_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_17_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_17_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_18_clock; // @[pe.scala 184:13]
  wire  PE_18_reset; // @[pe.scala 184:13]
  wire  PE_18_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_18_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_18_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_18_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_18_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_18_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_18_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_18_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_18_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_18_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_18_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_18_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_18_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_18_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_18_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_19_clock; // @[pe.scala 184:13]
  wire  PE_19_reset; // @[pe.scala 184:13]
  wire  PE_19_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_19_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_19_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_19_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_19_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_19_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_19_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_19_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_19_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_19_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_19_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_19_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_19_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_19_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_19_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_20_clock; // @[pe.scala 184:13]
  wire  PE_20_reset; // @[pe.scala 184:13]
  wire  PE_20_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_20_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_20_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_20_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_20_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_20_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_20_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_20_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_20_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_20_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_20_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_20_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_20_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_20_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_20_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_21_clock; // @[pe.scala 184:13]
  wire  PE_21_reset; // @[pe.scala 184:13]
  wire  PE_21_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_21_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_21_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_21_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_21_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_21_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_21_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_21_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_21_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_21_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_21_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_21_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_21_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_21_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_21_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_22_clock; // @[pe.scala 184:13]
  wire  PE_22_reset; // @[pe.scala 184:13]
  wire  PE_22_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_22_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_22_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_22_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_22_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_22_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_22_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_22_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_22_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_22_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_22_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_22_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_22_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_22_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_22_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_23_clock; // @[pe.scala 184:13]
  wire  PE_23_reset; // @[pe.scala 184:13]
  wire  PE_23_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_23_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_23_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_23_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_23_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_23_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_23_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_23_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_23_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_23_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_23_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_23_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_23_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_23_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_23_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_24_clock; // @[pe.scala 184:13]
  wire  PE_24_reset; // @[pe.scala 184:13]
  wire  PE_24_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_24_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_24_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_24_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_24_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_24_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_24_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_24_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_24_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_24_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_24_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_24_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_24_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_24_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_24_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_25_clock; // @[pe.scala 184:13]
  wire  PE_25_reset; // @[pe.scala 184:13]
  wire  PE_25_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_25_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_25_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_25_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_25_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_25_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_25_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_25_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_25_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_25_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_25_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_25_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_25_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_25_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_25_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_26_clock; // @[pe.scala 184:13]
  wire  PE_26_reset; // @[pe.scala 184:13]
  wire  PE_26_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_26_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_26_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_26_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_26_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_26_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_26_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_26_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_26_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_26_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_26_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_26_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_26_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_26_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_26_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_27_clock; // @[pe.scala 184:13]
  wire  PE_27_reset; // @[pe.scala 184:13]
  wire  PE_27_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_27_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_27_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_27_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_27_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_27_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_27_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_27_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_27_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_27_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_27_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_27_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_27_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_27_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_27_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_28_clock; // @[pe.scala 184:13]
  wire  PE_28_reset; // @[pe.scala 184:13]
  wire  PE_28_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_28_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_28_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_28_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_28_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_28_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_28_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_28_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_28_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_28_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_28_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_28_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_28_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_28_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_28_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_29_clock; // @[pe.scala 184:13]
  wire  PE_29_reset; // @[pe.scala 184:13]
  wire  PE_29_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_29_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_29_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_29_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_29_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_29_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_29_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_29_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_29_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_29_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_29_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_29_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_29_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_29_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_29_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_30_clock; // @[pe.scala 184:13]
  wire  PE_30_reset; // @[pe.scala 184:13]
  wire  PE_30_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_30_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_30_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_30_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_30_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_30_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_30_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_30_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_30_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_30_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_30_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_30_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_30_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_30_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_30_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_31_clock; // @[pe.scala 184:13]
  wire  PE_31_reset; // @[pe.scala 184:13]
  wire  PE_31_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_31_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_31_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_31_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_31_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_31_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_31_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_31_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_31_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_31_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_31_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_31_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_31_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_31_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_31_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_32_clock; // @[pe.scala 184:13]
  wire  PE_32_reset; // @[pe.scala 184:13]
  wire  PE_32_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_32_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_32_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_32_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_32_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_32_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_32_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_32_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_32_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_32_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_32_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_32_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_32_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_32_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_32_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_33_clock; // @[pe.scala 184:13]
  wire  PE_33_reset; // @[pe.scala 184:13]
  wire  PE_33_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_33_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_33_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_33_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_33_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_33_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_33_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_33_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_33_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_33_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_33_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_33_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_33_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_33_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_33_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_34_clock; // @[pe.scala 184:13]
  wire  PE_34_reset; // @[pe.scala 184:13]
  wire  PE_34_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_34_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_34_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_34_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_34_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_34_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_34_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_34_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_34_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_34_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_34_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_34_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_34_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_34_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_34_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_35_clock; // @[pe.scala 184:13]
  wire  PE_35_reset; // @[pe.scala 184:13]
  wire  PE_35_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_35_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_35_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_35_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_35_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_35_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_35_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_35_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_35_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_35_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_35_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_35_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_35_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_35_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_35_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_36_clock; // @[pe.scala 184:13]
  wire  PE_36_reset; // @[pe.scala 184:13]
  wire  PE_36_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_36_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_36_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_36_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_36_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_36_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_36_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_36_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_36_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_36_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_36_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_36_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_36_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_36_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_36_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_37_clock; // @[pe.scala 184:13]
  wire  PE_37_reset; // @[pe.scala 184:13]
  wire  PE_37_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_37_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_37_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_37_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_37_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_37_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_37_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_37_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_37_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_37_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_37_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_37_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_37_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_37_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_37_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_38_clock; // @[pe.scala 184:13]
  wire  PE_38_reset; // @[pe.scala 184:13]
  wire  PE_38_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_38_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_38_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_38_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_38_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_38_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_38_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_38_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_38_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_38_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_38_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_38_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_38_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_38_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_38_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_39_clock; // @[pe.scala 184:13]
  wire  PE_39_reset; // @[pe.scala 184:13]
  wire  PE_39_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_39_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_39_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_39_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_39_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_39_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_39_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_39_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_39_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_39_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_39_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_39_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_39_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_39_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_39_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_40_clock; // @[pe.scala 184:13]
  wire  PE_40_reset; // @[pe.scala 184:13]
  wire  PE_40_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_40_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_40_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_40_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_40_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_40_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_40_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_40_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_40_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_40_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_40_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_40_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_40_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_40_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_40_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_41_clock; // @[pe.scala 184:13]
  wire  PE_41_reset; // @[pe.scala 184:13]
  wire  PE_41_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_41_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_41_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_41_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_41_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_41_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_41_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_41_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_41_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_41_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_41_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_41_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_41_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_41_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_41_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_42_clock; // @[pe.scala 184:13]
  wire  PE_42_reset; // @[pe.scala 184:13]
  wire  PE_42_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_42_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_42_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_42_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_42_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_42_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_42_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_42_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_42_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_42_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_42_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_42_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_42_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_42_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_42_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_43_clock; // @[pe.scala 184:13]
  wire  PE_43_reset; // @[pe.scala 184:13]
  wire  PE_43_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_43_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_43_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_43_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_43_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_43_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_43_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_43_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_43_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_43_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_43_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_43_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_43_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_43_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_43_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_44_clock; // @[pe.scala 184:13]
  wire  PE_44_reset; // @[pe.scala 184:13]
  wire  PE_44_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_44_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_44_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_44_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_44_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_44_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_44_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_44_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_44_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_44_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_44_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_44_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_44_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_44_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_44_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_45_clock; // @[pe.scala 184:13]
  wire  PE_45_reset; // @[pe.scala 184:13]
  wire  PE_45_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_45_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_45_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_45_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_45_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_45_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_45_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_45_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_45_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_45_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_45_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_45_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_45_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_45_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_45_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_46_clock; // @[pe.scala 184:13]
  wire  PE_46_reset; // @[pe.scala 184:13]
  wire  PE_46_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_46_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_46_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_46_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_46_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_46_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_46_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_46_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_46_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_46_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_46_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_46_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_46_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_46_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_46_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_47_clock; // @[pe.scala 184:13]
  wire  PE_47_reset; // @[pe.scala 184:13]
  wire  PE_47_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_47_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_47_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_47_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_47_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_47_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_47_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_47_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_47_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_47_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_47_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_47_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_47_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_47_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_47_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_48_clock; // @[pe.scala 184:13]
  wire  PE_48_reset; // @[pe.scala 184:13]
  wire  PE_48_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_48_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_48_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_48_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_48_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_48_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_48_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_48_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_48_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_48_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_48_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_48_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_48_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_48_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_48_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_49_clock; // @[pe.scala 184:13]
  wire  PE_49_reset; // @[pe.scala 184:13]
  wire  PE_49_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_49_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_49_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_49_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_49_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_49_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_49_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_49_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_49_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_49_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_49_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_49_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_49_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_49_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_49_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_50_clock; // @[pe.scala 184:13]
  wire  PE_50_reset; // @[pe.scala 184:13]
  wire  PE_50_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_50_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_50_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_50_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_50_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_50_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_50_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_50_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_50_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_50_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_50_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_50_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_50_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_50_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_50_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_51_clock; // @[pe.scala 184:13]
  wire  PE_51_reset; // @[pe.scala 184:13]
  wire  PE_51_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_51_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_51_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_51_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_51_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_51_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_51_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_51_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_51_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_51_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_51_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_51_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_51_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_51_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_51_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_52_clock; // @[pe.scala 184:13]
  wire  PE_52_reset; // @[pe.scala 184:13]
  wire  PE_52_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_52_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_52_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_52_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_52_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_52_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_52_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_52_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_52_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_52_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_52_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_52_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_52_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_52_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_52_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_53_clock; // @[pe.scala 184:13]
  wire  PE_53_reset; // @[pe.scala 184:13]
  wire  PE_53_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_53_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_53_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_53_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_53_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_53_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_53_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_53_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_53_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_53_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_53_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_53_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_53_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_53_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_53_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_54_clock; // @[pe.scala 184:13]
  wire  PE_54_reset; // @[pe.scala 184:13]
  wire  PE_54_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_54_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_54_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_54_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_54_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_54_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_54_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_54_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_54_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_54_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_54_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_54_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_54_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_54_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_54_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_55_clock; // @[pe.scala 184:13]
  wire  PE_55_reset; // @[pe.scala 184:13]
  wire  PE_55_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_55_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_55_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_55_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_55_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_55_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_55_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_55_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_55_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_55_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_55_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_55_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_55_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_55_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_55_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_56_clock; // @[pe.scala 184:13]
  wire  PE_56_reset; // @[pe.scala 184:13]
  wire  PE_56_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_56_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_56_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_56_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_56_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_56_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_56_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_56_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_56_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_56_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_56_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_56_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_56_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_56_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_56_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_57_clock; // @[pe.scala 184:13]
  wire  PE_57_reset; // @[pe.scala 184:13]
  wire  PE_57_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_57_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_57_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_57_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_57_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_57_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_57_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_57_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_57_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_57_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_57_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_57_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_57_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_57_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_57_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_58_clock; // @[pe.scala 184:13]
  wire  PE_58_reset; // @[pe.scala 184:13]
  wire  PE_58_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_58_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_58_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_58_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_58_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_58_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_58_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_58_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_58_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_58_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_58_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_58_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_58_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_58_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_58_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_59_clock; // @[pe.scala 184:13]
  wire  PE_59_reset; // @[pe.scala 184:13]
  wire  PE_59_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_59_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_59_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_59_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_59_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_59_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_59_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_59_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_59_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_59_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_59_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_59_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_59_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_59_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_59_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_60_clock; // @[pe.scala 184:13]
  wire  PE_60_reset; // @[pe.scala 184:13]
  wire  PE_60_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_60_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_60_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_60_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_60_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_60_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_60_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_60_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_60_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_60_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_60_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_60_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_60_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_60_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_60_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_61_clock; // @[pe.scala 184:13]
  wire  PE_61_reset; // @[pe.scala 184:13]
  wire  PE_61_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_61_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_61_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_61_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_61_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_61_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_61_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_61_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_61_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_61_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_61_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_61_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_61_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_61_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_61_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_62_clock; // @[pe.scala 184:13]
  wire  PE_62_reset; // @[pe.scala 184:13]
  wire  PE_62_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_62_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_62_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_62_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_62_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_62_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_62_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_62_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_62_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_62_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_62_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_62_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_62_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_62_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_62_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_63_clock; // @[pe.scala 184:13]
  wire  PE_63_reset; // @[pe.scala 184:13]
  wire  PE_63_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_63_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_63_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_63_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_63_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_63_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_63_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_63_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_63_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_63_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_63_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_63_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_63_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_63_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_63_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_64_clock; // @[pe.scala 184:13]
  wire  PE_64_reset; // @[pe.scala 184:13]
  wire  PE_64_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_64_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_64_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_64_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_64_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_64_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_64_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_64_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_64_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_64_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_64_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_64_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_64_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_64_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_64_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_65_clock; // @[pe.scala 184:13]
  wire  PE_65_reset; // @[pe.scala 184:13]
  wire  PE_65_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_65_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_65_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_65_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_65_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_65_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_65_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_65_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_65_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_65_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_65_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_65_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_65_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_65_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_65_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_66_clock; // @[pe.scala 184:13]
  wire  PE_66_reset; // @[pe.scala 184:13]
  wire  PE_66_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_66_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_66_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_66_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_66_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_66_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_66_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_66_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_66_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_66_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_66_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_66_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_66_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_66_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_66_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_67_clock; // @[pe.scala 184:13]
  wire  PE_67_reset; // @[pe.scala 184:13]
  wire  PE_67_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_67_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_67_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_67_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_67_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_67_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_67_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_67_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_67_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_67_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_67_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_67_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_67_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_67_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_67_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_68_clock; // @[pe.scala 184:13]
  wire  PE_68_reset; // @[pe.scala 184:13]
  wire  PE_68_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_68_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_68_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_68_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_68_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_68_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_68_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_68_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_68_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_68_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_68_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_68_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_68_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_68_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_68_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_69_clock; // @[pe.scala 184:13]
  wire  PE_69_reset; // @[pe.scala 184:13]
  wire  PE_69_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_69_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_69_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_69_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_69_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_69_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_69_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_69_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_69_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_69_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_69_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_69_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_69_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_69_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_69_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_70_clock; // @[pe.scala 184:13]
  wire  PE_70_reset; // @[pe.scala 184:13]
  wire  PE_70_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_70_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_70_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_70_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_70_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_70_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_70_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_70_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_70_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_70_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_70_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_70_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_70_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_70_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_70_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_71_clock; // @[pe.scala 184:13]
  wire  PE_71_reset; // @[pe.scala 184:13]
  wire  PE_71_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_71_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_71_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_71_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_71_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_71_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_71_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_71_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_71_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_71_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_71_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_71_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_71_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_71_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_71_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_72_clock; // @[pe.scala 184:13]
  wire  PE_72_reset; // @[pe.scala 184:13]
  wire  PE_72_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_72_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_72_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_72_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_72_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_72_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_72_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_72_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_72_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_72_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_72_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_72_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_72_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_72_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_72_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_73_clock; // @[pe.scala 184:13]
  wire  PE_73_reset; // @[pe.scala 184:13]
  wire  PE_73_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_73_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_73_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_73_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_73_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_73_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_73_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_73_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_73_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_73_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_73_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_73_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_73_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_73_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_73_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_74_clock; // @[pe.scala 184:13]
  wire  PE_74_reset; // @[pe.scala 184:13]
  wire  PE_74_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_74_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_74_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_74_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_74_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_74_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_74_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_74_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_74_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_74_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_74_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_74_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_74_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_74_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_74_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_75_clock; // @[pe.scala 184:13]
  wire  PE_75_reset; // @[pe.scala 184:13]
  wire  PE_75_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_75_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_75_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_75_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_75_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_75_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_75_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_75_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_75_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_75_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_75_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_75_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_75_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_75_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_75_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_76_clock; // @[pe.scala 184:13]
  wire  PE_76_reset; // @[pe.scala 184:13]
  wire  PE_76_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_76_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_76_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_76_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_76_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_76_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_76_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_76_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_76_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_76_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_76_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_76_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_76_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_76_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_76_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_77_clock; // @[pe.scala 184:13]
  wire  PE_77_reset; // @[pe.scala 184:13]
  wire  PE_77_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_77_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_77_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_77_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_77_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_77_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_77_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_77_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_77_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_77_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_77_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_77_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_77_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_77_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_77_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_78_clock; // @[pe.scala 184:13]
  wire  PE_78_reset; // @[pe.scala 184:13]
  wire  PE_78_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_78_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_78_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_78_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_78_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_78_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_78_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_78_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_78_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_78_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_78_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_78_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_78_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_78_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_78_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_79_clock; // @[pe.scala 184:13]
  wire  PE_79_reset; // @[pe.scala 184:13]
  wire  PE_79_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_79_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_79_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_79_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_79_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_79_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_79_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_79_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_79_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_79_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_79_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_79_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_79_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_79_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_79_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_80_clock; // @[pe.scala 184:13]
  wire  PE_80_reset; // @[pe.scala 184:13]
  wire  PE_80_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_80_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_80_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_80_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_80_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_80_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_80_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_80_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_80_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_80_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_80_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_80_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_80_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_80_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_80_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_81_clock; // @[pe.scala 184:13]
  wire  PE_81_reset; // @[pe.scala 184:13]
  wire  PE_81_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_81_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_81_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_81_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_81_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_81_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_81_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_81_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_81_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_81_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_81_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_81_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_81_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_81_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_81_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_82_clock; // @[pe.scala 184:13]
  wire  PE_82_reset; // @[pe.scala 184:13]
  wire  PE_82_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_82_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_82_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_82_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_82_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_82_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_82_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_82_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_82_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_82_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_82_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_82_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_82_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_82_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_82_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_83_clock; // @[pe.scala 184:13]
  wire  PE_83_reset; // @[pe.scala 184:13]
  wire  PE_83_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_83_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_83_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_83_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_83_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_83_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_83_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_83_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_83_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_83_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_83_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_83_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_83_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_83_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_83_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_84_clock; // @[pe.scala 184:13]
  wire  PE_84_reset; // @[pe.scala 184:13]
  wire  PE_84_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_84_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_84_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_84_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_84_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_84_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_84_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_84_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_84_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_84_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_84_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_84_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_84_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_84_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_84_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_85_clock; // @[pe.scala 184:13]
  wire  PE_85_reset; // @[pe.scala 184:13]
  wire  PE_85_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_85_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_85_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_85_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_85_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_85_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_85_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_85_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_85_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_85_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_85_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_85_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_85_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_85_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_85_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_86_clock; // @[pe.scala 184:13]
  wire  PE_86_reset; // @[pe.scala 184:13]
  wire  PE_86_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_86_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_86_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_86_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_86_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_86_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_86_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_86_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_86_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_86_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_86_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_86_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_86_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_86_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_86_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_87_clock; // @[pe.scala 184:13]
  wire  PE_87_reset; // @[pe.scala 184:13]
  wire  PE_87_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_87_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_87_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_87_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_87_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_87_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_87_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_87_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_87_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_87_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_87_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_87_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_87_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_87_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_87_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_88_clock; // @[pe.scala 184:13]
  wire  PE_88_reset; // @[pe.scala 184:13]
  wire  PE_88_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_88_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_88_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_88_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_88_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_88_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_88_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_88_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_88_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_88_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_88_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_88_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_88_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_88_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_88_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_89_clock; // @[pe.scala 184:13]
  wire  PE_89_reset; // @[pe.scala 184:13]
  wire  PE_89_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_89_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_89_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_89_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_89_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_89_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_89_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_89_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_89_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_89_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_89_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_89_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_89_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_89_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_89_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_90_clock; // @[pe.scala 184:13]
  wire  PE_90_reset; // @[pe.scala 184:13]
  wire  PE_90_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_90_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_90_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_90_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_90_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_90_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_90_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_90_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_90_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_90_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_90_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_90_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_90_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_90_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_90_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_91_clock; // @[pe.scala 184:13]
  wire  PE_91_reset; // @[pe.scala 184:13]
  wire  PE_91_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_91_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_91_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_91_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_91_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_91_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_91_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_91_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_91_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_91_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_91_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_91_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_91_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_91_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_91_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_92_clock; // @[pe.scala 184:13]
  wire  PE_92_reset; // @[pe.scala 184:13]
  wire  PE_92_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_92_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_92_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_92_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_92_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_92_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_92_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_92_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_92_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_92_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_92_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_92_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_92_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_92_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_92_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_93_clock; // @[pe.scala 184:13]
  wire  PE_93_reset; // @[pe.scala 184:13]
  wire  PE_93_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_93_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_93_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_93_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_93_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_93_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_93_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_93_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_93_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_93_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_93_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_93_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_93_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_93_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_93_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_94_clock; // @[pe.scala 184:13]
  wire  PE_94_reset; // @[pe.scala 184:13]
  wire  PE_94_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_94_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_94_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_94_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_94_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_94_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_94_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_94_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_94_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_94_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_94_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_94_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_94_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_94_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_94_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_95_clock; // @[pe.scala 184:13]
  wire  PE_95_reset; // @[pe.scala 184:13]
  wire  PE_95_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_95_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_95_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_95_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_95_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_95_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_95_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_95_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_95_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_95_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_95_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_95_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_95_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_95_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_95_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_96_clock; // @[pe.scala 184:13]
  wire  PE_96_reset; // @[pe.scala 184:13]
  wire  PE_96_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_96_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_96_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_96_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_96_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_96_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_96_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_96_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_96_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_96_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_96_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_96_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_96_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_96_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_96_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_97_clock; // @[pe.scala 184:13]
  wire  PE_97_reset; // @[pe.scala 184:13]
  wire  PE_97_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_97_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_97_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_97_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_97_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_97_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_97_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_97_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_97_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_97_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_97_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_97_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_97_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_97_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_97_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_98_clock; // @[pe.scala 184:13]
  wire  PE_98_reset; // @[pe.scala 184:13]
  wire  PE_98_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_98_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_98_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_98_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_98_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_98_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_98_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_98_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_98_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_98_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_98_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_98_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_98_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_98_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_98_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_99_clock; // @[pe.scala 184:13]
  wire  PE_99_reset; // @[pe.scala 184:13]
  wire  PE_99_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_99_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_99_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_99_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_99_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_99_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_99_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_99_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_99_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_99_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_99_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_99_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_99_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_99_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_99_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_100_clock; // @[pe.scala 184:13]
  wire  PE_100_reset; // @[pe.scala 184:13]
  wire  PE_100_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_100_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_100_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_100_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_100_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_100_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_100_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_100_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_100_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_100_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_100_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_100_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_100_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_100_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_100_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_101_clock; // @[pe.scala 184:13]
  wire  PE_101_reset; // @[pe.scala 184:13]
  wire  PE_101_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_101_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_101_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_101_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_101_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_101_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_101_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_101_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_101_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_101_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_101_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_101_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_101_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_101_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_101_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_102_clock; // @[pe.scala 184:13]
  wire  PE_102_reset; // @[pe.scala 184:13]
  wire  PE_102_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_102_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_102_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_102_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_102_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_102_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_102_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_102_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_102_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_102_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_102_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_102_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_102_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_102_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_102_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_103_clock; // @[pe.scala 184:13]
  wire  PE_103_reset; // @[pe.scala 184:13]
  wire  PE_103_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_103_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_103_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_103_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_103_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_103_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_103_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_103_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_103_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_103_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_103_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_103_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_103_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_103_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_103_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_104_clock; // @[pe.scala 184:13]
  wire  PE_104_reset; // @[pe.scala 184:13]
  wire  PE_104_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_104_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_104_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_104_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_104_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_104_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_104_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_104_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_104_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_104_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_104_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_104_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_104_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_104_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_104_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_105_clock; // @[pe.scala 184:13]
  wire  PE_105_reset; // @[pe.scala 184:13]
  wire  PE_105_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_105_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_105_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_105_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_105_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_105_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_105_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_105_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_105_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_105_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_105_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_105_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_105_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_105_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_105_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_106_clock; // @[pe.scala 184:13]
  wire  PE_106_reset; // @[pe.scala 184:13]
  wire  PE_106_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_106_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_106_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_106_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_106_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_106_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_106_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_106_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_106_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_106_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_106_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_106_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_106_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_106_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_106_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_107_clock; // @[pe.scala 184:13]
  wire  PE_107_reset; // @[pe.scala 184:13]
  wire  PE_107_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_107_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_107_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_107_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_107_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_107_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_107_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_107_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_107_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_107_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_107_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_107_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_107_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_107_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_107_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_108_clock; // @[pe.scala 184:13]
  wire  PE_108_reset; // @[pe.scala 184:13]
  wire  PE_108_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_108_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_108_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_108_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_108_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_108_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_108_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_108_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_108_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_108_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_108_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_108_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_108_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_108_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_108_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_109_clock; // @[pe.scala 184:13]
  wire  PE_109_reset; // @[pe.scala 184:13]
  wire  PE_109_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_109_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_109_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_109_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_109_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_109_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_109_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_109_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_109_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_109_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_109_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_109_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_109_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_109_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_109_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_110_clock; // @[pe.scala 184:13]
  wire  PE_110_reset; // @[pe.scala 184:13]
  wire  PE_110_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_110_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_110_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_110_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_110_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_110_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_110_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_110_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_110_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_110_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_110_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_110_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_110_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_110_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_110_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_111_clock; // @[pe.scala 184:13]
  wire  PE_111_reset; // @[pe.scala 184:13]
  wire  PE_111_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_111_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_111_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_111_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_111_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_111_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_111_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_111_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_111_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_111_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_111_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_111_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_111_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_111_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_111_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_112_clock; // @[pe.scala 184:13]
  wire  PE_112_reset; // @[pe.scala 184:13]
  wire  PE_112_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_112_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_112_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_112_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_112_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_112_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_112_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_112_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_112_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_112_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_112_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_112_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_112_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_112_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_112_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_113_clock; // @[pe.scala 184:13]
  wire  PE_113_reset; // @[pe.scala 184:13]
  wire  PE_113_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_113_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_113_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_113_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_113_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_113_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_113_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_113_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_113_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_113_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_113_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_113_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_113_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_113_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_113_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_114_clock; // @[pe.scala 184:13]
  wire  PE_114_reset; // @[pe.scala 184:13]
  wire  PE_114_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_114_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_114_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_114_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_114_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_114_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_114_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_114_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_114_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_114_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_114_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_114_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_114_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_114_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_114_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_115_clock; // @[pe.scala 184:13]
  wire  PE_115_reset; // @[pe.scala 184:13]
  wire  PE_115_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_115_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_115_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_115_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_115_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_115_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_115_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_115_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_115_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_115_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_115_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_115_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_115_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_115_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_115_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_116_clock; // @[pe.scala 184:13]
  wire  PE_116_reset; // @[pe.scala 184:13]
  wire  PE_116_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_116_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_116_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_116_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_116_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_116_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_116_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_116_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_116_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_116_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_116_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_116_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_116_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_116_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_116_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_117_clock; // @[pe.scala 184:13]
  wire  PE_117_reset; // @[pe.scala 184:13]
  wire  PE_117_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_117_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_117_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_117_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_117_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_117_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_117_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_117_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_117_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_117_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_117_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_117_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_117_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_117_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_117_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_118_clock; // @[pe.scala 184:13]
  wire  PE_118_reset; // @[pe.scala 184:13]
  wire  PE_118_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_118_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_118_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_118_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_118_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_118_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_118_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_118_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_118_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_118_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_118_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_118_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_118_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_118_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_118_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_119_clock; // @[pe.scala 184:13]
  wire  PE_119_reset; // @[pe.scala 184:13]
  wire  PE_119_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_119_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_119_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_119_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_119_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_119_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_119_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_119_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_119_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_119_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_119_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_119_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_119_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_119_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_119_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_120_clock; // @[pe.scala 184:13]
  wire  PE_120_reset; // @[pe.scala 184:13]
  wire  PE_120_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_120_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_120_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_120_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_120_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_120_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_120_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_120_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_120_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_120_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_120_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_120_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_120_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_120_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_120_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_121_clock; // @[pe.scala 184:13]
  wire  PE_121_reset; // @[pe.scala 184:13]
  wire  PE_121_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_121_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_121_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_121_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_121_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_121_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_121_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_121_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_121_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_121_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_121_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_121_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_121_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_121_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_121_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_122_clock; // @[pe.scala 184:13]
  wire  PE_122_reset; // @[pe.scala 184:13]
  wire  PE_122_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_122_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_122_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_122_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_122_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_122_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_122_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_122_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_122_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_122_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_122_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_122_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_122_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_122_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_122_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_123_clock; // @[pe.scala 184:13]
  wire  PE_123_reset; // @[pe.scala 184:13]
  wire  PE_123_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_123_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_123_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_123_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_123_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_123_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_123_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_123_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_123_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_123_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_123_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_123_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_123_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_123_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_123_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_124_clock; // @[pe.scala 184:13]
  wire  PE_124_reset; // @[pe.scala 184:13]
  wire  PE_124_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_124_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_124_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_124_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_124_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_124_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_124_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_124_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_124_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_124_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_124_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_124_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_124_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_124_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_124_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_125_clock; // @[pe.scala 184:13]
  wire  PE_125_reset; // @[pe.scala 184:13]
  wire  PE_125_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_125_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_125_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_125_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_125_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_125_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_125_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_125_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_125_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_125_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_125_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_125_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_125_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_125_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_125_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_126_clock; // @[pe.scala 184:13]
  wire  PE_126_reset; // @[pe.scala 184:13]
  wire  PE_126_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_126_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_126_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_126_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_126_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_126_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_126_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_126_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_126_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_126_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_126_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_126_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_126_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_126_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_126_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_127_clock; // @[pe.scala 184:13]
  wire  PE_127_reset; // @[pe.scala 184:13]
  wire  PE_127_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_127_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_127_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_127_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_127_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_127_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_127_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_127_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_127_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_127_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_127_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_127_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_127_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_127_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_127_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_128_clock; // @[pe.scala 184:13]
  wire  PE_128_reset; // @[pe.scala 184:13]
  wire  PE_128_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_128_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_128_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_128_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_128_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_128_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_128_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_128_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_128_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_128_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_128_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_128_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_128_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_128_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_128_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_129_clock; // @[pe.scala 184:13]
  wire  PE_129_reset; // @[pe.scala 184:13]
  wire  PE_129_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_129_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_129_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_129_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_129_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_129_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_129_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_129_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_129_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_129_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_129_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_129_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_129_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_129_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_129_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_130_clock; // @[pe.scala 184:13]
  wire  PE_130_reset; // @[pe.scala 184:13]
  wire  PE_130_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_130_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_130_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_130_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_130_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_130_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_130_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_130_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_130_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_130_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_130_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_130_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_130_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_130_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_130_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_131_clock; // @[pe.scala 184:13]
  wire  PE_131_reset; // @[pe.scala 184:13]
  wire  PE_131_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_131_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_131_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_131_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_131_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_131_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_131_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_131_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_131_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_131_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_131_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_131_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_131_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_131_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_131_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_132_clock; // @[pe.scala 184:13]
  wire  PE_132_reset; // @[pe.scala 184:13]
  wire  PE_132_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_132_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_132_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_132_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_132_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_132_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_132_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_132_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_132_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_132_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_132_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_132_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_132_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_132_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_132_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_133_clock; // @[pe.scala 184:13]
  wire  PE_133_reset; // @[pe.scala 184:13]
  wire  PE_133_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_133_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_133_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_133_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_133_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_133_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_133_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_133_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_133_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_133_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_133_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_133_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_133_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_133_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_133_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_134_clock; // @[pe.scala 184:13]
  wire  PE_134_reset; // @[pe.scala 184:13]
  wire  PE_134_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_134_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_134_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_134_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_134_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_134_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_134_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_134_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_134_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_134_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_134_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_134_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_134_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_134_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_134_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_135_clock; // @[pe.scala 184:13]
  wire  PE_135_reset; // @[pe.scala 184:13]
  wire  PE_135_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_135_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_135_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_135_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_135_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_135_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_135_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_135_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_135_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_135_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_135_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_135_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_135_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_135_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_135_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_136_clock; // @[pe.scala 184:13]
  wire  PE_136_reset; // @[pe.scala 184:13]
  wire  PE_136_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_136_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_136_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_136_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_136_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_136_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_136_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_136_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_136_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_136_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_136_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_136_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_136_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_136_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_136_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_137_clock; // @[pe.scala 184:13]
  wire  PE_137_reset; // @[pe.scala 184:13]
  wire  PE_137_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_137_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_137_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_137_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_137_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_137_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_137_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_137_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_137_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_137_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_137_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_137_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_137_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_137_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_137_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_138_clock; // @[pe.scala 184:13]
  wire  PE_138_reset; // @[pe.scala 184:13]
  wire  PE_138_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_138_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_138_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_138_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_138_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_138_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_138_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_138_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_138_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_138_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_138_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_138_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_138_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_138_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_138_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_139_clock; // @[pe.scala 184:13]
  wire  PE_139_reset; // @[pe.scala 184:13]
  wire  PE_139_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_139_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_139_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_139_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_139_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_139_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_139_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_139_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_139_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_139_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_139_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_139_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_139_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_139_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_139_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_140_clock; // @[pe.scala 184:13]
  wire  PE_140_reset; // @[pe.scala 184:13]
  wire  PE_140_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_140_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_140_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_140_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_140_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_140_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_140_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_140_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_140_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_140_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_140_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_140_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_140_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_140_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_140_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_141_clock; // @[pe.scala 184:13]
  wire  PE_141_reset; // @[pe.scala 184:13]
  wire  PE_141_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_141_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_141_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_141_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_141_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_141_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_141_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_141_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_141_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_141_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_141_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_141_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_141_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_141_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_141_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_142_clock; // @[pe.scala 184:13]
  wire  PE_142_reset; // @[pe.scala 184:13]
  wire  PE_142_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_142_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_142_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_142_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_142_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_142_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_142_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_142_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_142_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_142_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_142_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_142_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_142_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_142_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_142_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_143_clock; // @[pe.scala 184:13]
  wire  PE_143_reset; // @[pe.scala 184:13]
  wire  PE_143_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_143_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_143_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_143_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_143_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_143_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_143_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_143_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_143_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_143_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_143_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_143_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_143_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_143_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_143_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_144_clock; // @[pe.scala 184:13]
  wire  PE_144_reset; // @[pe.scala 184:13]
  wire  PE_144_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_144_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_144_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_144_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_144_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_144_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_144_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_144_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_144_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_144_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_144_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_144_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_144_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_144_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_144_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_145_clock; // @[pe.scala 184:13]
  wire  PE_145_reset; // @[pe.scala 184:13]
  wire  PE_145_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_145_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_145_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_145_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_145_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_145_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_145_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_145_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_145_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_145_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_145_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_145_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_145_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_145_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_145_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_146_clock; // @[pe.scala 184:13]
  wire  PE_146_reset; // @[pe.scala 184:13]
  wire  PE_146_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_146_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_146_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_146_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_146_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_146_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_146_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_146_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_146_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_146_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_146_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_146_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_146_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_146_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_146_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_147_clock; // @[pe.scala 184:13]
  wire  PE_147_reset; // @[pe.scala 184:13]
  wire  PE_147_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_147_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_147_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_147_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_147_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_147_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_147_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_147_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_147_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_147_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_147_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_147_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_147_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_147_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_147_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_148_clock; // @[pe.scala 184:13]
  wire  PE_148_reset; // @[pe.scala 184:13]
  wire  PE_148_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_148_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_148_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_148_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_148_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_148_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_148_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_148_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_148_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_148_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_148_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_148_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_148_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_148_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_148_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_149_clock; // @[pe.scala 184:13]
  wire  PE_149_reset; // @[pe.scala 184:13]
  wire  PE_149_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_149_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_149_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_149_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_149_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_149_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_149_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_149_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_149_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_149_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_149_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_149_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_149_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_149_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_149_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_150_clock; // @[pe.scala 184:13]
  wire  PE_150_reset; // @[pe.scala 184:13]
  wire  PE_150_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_150_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_150_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_150_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_150_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_150_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_150_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_150_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_150_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_150_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_150_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_150_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_150_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_150_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_150_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_151_clock; // @[pe.scala 184:13]
  wire  PE_151_reset; // @[pe.scala 184:13]
  wire  PE_151_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_151_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_151_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_151_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_151_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_151_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_151_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_151_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_151_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_151_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_151_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_151_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_151_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_151_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_151_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_152_clock; // @[pe.scala 184:13]
  wire  PE_152_reset; // @[pe.scala 184:13]
  wire  PE_152_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_152_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_152_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_152_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_152_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_152_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_152_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_152_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_152_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_152_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_152_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_152_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_152_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_152_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_152_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_153_clock; // @[pe.scala 184:13]
  wire  PE_153_reset; // @[pe.scala 184:13]
  wire  PE_153_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_153_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_153_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_153_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_153_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_153_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_153_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_153_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_153_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_153_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_153_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_153_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_153_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_153_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_153_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_154_clock; // @[pe.scala 184:13]
  wire  PE_154_reset; // @[pe.scala 184:13]
  wire  PE_154_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_154_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_154_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_154_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_154_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_154_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_154_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_154_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_154_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_154_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_154_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_154_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_154_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_154_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_154_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_155_clock; // @[pe.scala 184:13]
  wire  PE_155_reset; // @[pe.scala 184:13]
  wire  PE_155_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_155_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_155_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_155_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_155_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_155_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_155_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_155_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_155_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_155_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_155_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_155_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_155_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_155_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_155_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_156_clock; // @[pe.scala 184:13]
  wire  PE_156_reset; // @[pe.scala 184:13]
  wire  PE_156_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_156_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_156_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_156_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_156_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_156_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_156_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_156_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_156_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_156_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_156_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_156_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_156_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_156_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_156_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_157_clock; // @[pe.scala 184:13]
  wire  PE_157_reset; // @[pe.scala 184:13]
  wire  PE_157_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_157_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_157_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_157_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_157_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_157_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_157_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_157_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_157_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_157_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_157_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_157_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_157_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_157_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_157_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_158_clock; // @[pe.scala 184:13]
  wire  PE_158_reset; // @[pe.scala 184:13]
  wire  PE_158_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_158_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_158_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_158_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_158_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_158_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_158_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_158_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_158_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_158_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_158_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_158_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_158_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_158_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_158_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_159_clock; // @[pe.scala 184:13]
  wire  PE_159_reset; // @[pe.scala 184:13]
  wire  PE_159_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_159_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_159_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_159_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_159_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_159_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_159_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_159_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_159_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_159_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_159_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_159_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_159_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_159_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_159_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_160_clock; // @[pe.scala 184:13]
  wire  PE_160_reset; // @[pe.scala 184:13]
  wire  PE_160_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_160_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_160_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_160_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_160_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_160_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_160_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_160_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_160_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_160_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_160_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_160_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_160_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_160_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_160_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_161_clock; // @[pe.scala 184:13]
  wire  PE_161_reset; // @[pe.scala 184:13]
  wire  PE_161_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_161_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_161_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_161_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_161_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_161_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_161_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_161_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_161_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_161_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_161_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_161_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_161_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_161_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_161_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_162_clock; // @[pe.scala 184:13]
  wire  PE_162_reset; // @[pe.scala 184:13]
  wire  PE_162_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_162_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_162_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_162_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_162_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_162_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_162_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_162_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_162_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_162_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_162_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_162_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_162_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_162_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_162_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_163_clock; // @[pe.scala 184:13]
  wire  PE_163_reset; // @[pe.scala 184:13]
  wire  PE_163_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_163_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_163_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_163_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_163_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_163_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_163_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_163_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_163_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_163_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_163_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_163_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_163_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_163_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_163_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PE_164_clock; // @[pe.scala 184:13]
  wire  PE_164_reset; // @[pe.scala 184:13]
  wire  PE_164_io_data_2_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_164_io_data_2_in_bits; // @[pe.scala 184:13]
  wire  PE_164_io_data_2_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_164_io_data_2_out_bits; // @[pe.scala 184:13]
  wire  PE_164_io_data_2_sig_stat2trans; // @[pe.scala 184:13]
  wire  PE_164_io_data_2_in_ready; // @[pe.scala 184:13]
  wire  PE_164_io_data_2_out_ready; // @[pe.scala 184:13]
  wire  PE_164_io_data_1_in_valid; // @[pe.scala 184:13]
  wire [255:0] PE_164_io_data_1_in_bits; // @[pe.scala 184:13]
  wire  PE_164_io_data_1_out_valid; // @[pe.scala 184:13]
  wire [255:0] PE_164_io_data_1_out_bits; // @[pe.scala 184:13]
  wire  PE_164_io_data_0_in_valid; // @[pe.scala 184:13]
  wire [31:0] PE_164_io_data_0_in_bits; // @[pe.scala 184:13]
  wire  PE_164_io_data_0_out_valid; // @[pe.scala 184:13]
  wire [31:0] PE_164_io_data_0_out_bits; // @[pe.scala 184:13]
  wire  PENetwork_io_to_pes_0_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_io_to_pes_0_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_io_to_pes_0_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_io_to_pes_0_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_io_to_pes_1_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_io_to_pes_1_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_io_to_pes_1_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_io_to_pes_1_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_io_to_pes_2_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_io_to_pes_2_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_io_to_pes_2_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_io_to_pes_2_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_io_to_pes_3_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_io_to_pes_3_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_io_to_pes_3_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_io_to_pes_3_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_io_to_pes_4_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_io_to_pes_4_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_io_to_pes_4_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_io_to_pes_4_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_io_to_pes_5_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_io_to_pes_5_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_io_to_pes_5_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_io_to_pes_5_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_io_to_pes_6_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_io_to_pes_6_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_io_to_pes_6_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_io_to_pes_6_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_io_to_pes_7_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_io_to_pes_7_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_io_to_pes_7_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_io_to_pes_7_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_io_to_pes_8_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_io_to_pes_8_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_io_to_pes_8_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_io_to_pes_8_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_io_to_pes_9_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_io_to_pes_9_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_io_to_pes_9_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_io_to_pes_9_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_io_to_pes_10_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_io_to_pes_10_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_io_to_pes_10_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_io_to_pes_10_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_io_to_pes_11_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_io_to_pes_11_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_io_to_pes_11_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_io_to_pes_11_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_io_to_pes_12_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_io_to_pes_12_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_io_to_pes_12_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_io_to_pes_12_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_io_to_pes_13_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_io_to_pes_13_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_io_to_pes_13_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_io_to_pes_13_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_io_to_pes_14_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_io_to_pes_14_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_io_to_mem_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_io_to_mem_bits; // @[pe.scala 227:13]
  wire  PENetwork_1_io_to_pes_0_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_1_io_to_pes_0_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_1_io_to_pes_0_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_1_io_to_pes_0_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_1_io_to_pes_1_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_1_io_to_pes_1_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_1_io_to_pes_1_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_1_io_to_pes_1_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_1_io_to_pes_2_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_1_io_to_pes_2_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_1_io_to_pes_2_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_1_io_to_pes_2_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_1_io_to_pes_3_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_1_io_to_pes_3_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_1_io_to_pes_3_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_1_io_to_pes_3_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_1_io_to_pes_4_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_1_io_to_pes_4_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_1_io_to_pes_4_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_1_io_to_pes_4_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_1_io_to_pes_5_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_1_io_to_pes_5_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_1_io_to_pes_5_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_1_io_to_pes_5_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_1_io_to_pes_6_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_1_io_to_pes_6_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_1_io_to_pes_6_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_1_io_to_pes_6_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_1_io_to_pes_7_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_1_io_to_pes_7_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_1_io_to_pes_7_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_1_io_to_pes_7_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_1_io_to_pes_8_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_1_io_to_pes_8_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_1_io_to_pes_8_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_1_io_to_pes_8_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_1_io_to_pes_9_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_1_io_to_pes_9_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_1_io_to_pes_9_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_1_io_to_pes_9_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_1_io_to_pes_10_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_1_io_to_pes_10_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_1_io_to_pes_10_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_1_io_to_pes_10_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_1_io_to_pes_11_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_1_io_to_pes_11_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_1_io_to_pes_11_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_1_io_to_pes_11_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_1_io_to_pes_12_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_1_io_to_pes_12_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_1_io_to_pes_12_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_1_io_to_pes_12_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_1_io_to_pes_13_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_1_io_to_pes_13_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_1_io_to_pes_13_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_1_io_to_pes_13_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_1_io_to_pes_14_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_1_io_to_pes_14_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_1_io_to_mem_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_1_io_to_mem_bits; // @[pe.scala 227:13]
  wire  PENetwork_2_io_to_pes_0_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_2_io_to_pes_0_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_2_io_to_pes_0_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_2_io_to_pes_0_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_2_io_to_pes_1_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_2_io_to_pes_1_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_2_io_to_pes_1_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_2_io_to_pes_1_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_2_io_to_pes_2_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_2_io_to_pes_2_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_2_io_to_pes_2_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_2_io_to_pes_2_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_2_io_to_pes_3_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_2_io_to_pes_3_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_2_io_to_pes_3_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_2_io_to_pes_3_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_2_io_to_pes_4_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_2_io_to_pes_4_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_2_io_to_pes_4_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_2_io_to_pes_4_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_2_io_to_pes_5_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_2_io_to_pes_5_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_2_io_to_pes_5_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_2_io_to_pes_5_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_2_io_to_pes_6_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_2_io_to_pes_6_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_2_io_to_pes_6_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_2_io_to_pes_6_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_2_io_to_pes_7_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_2_io_to_pes_7_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_2_io_to_pes_7_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_2_io_to_pes_7_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_2_io_to_pes_8_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_2_io_to_pes_8_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_2_io_to_pes_8_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_2_io_to_pes_8_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_2_io_to_pes_9_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_2_io_to_pes_9_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_2_io_to_pes_9_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_2_io_to_pes_9_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_2_io_to_pes_10_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_2_io_to_pes_10_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_2_io_to_pes_10_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_2_io_to_pes_10_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_2_io_to_pes_11_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_2_io_to_pes_11_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_2_io_to_pes_11_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_2_io_to_pes_11_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_2_io_to_pes_12_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_2_io_to_pes_12_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_2_io_to_pes_12_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_2_io_to_pes_12_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_2_io_to_pes_13_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_2_io_to_pes_13_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_2_io_to_pes_13_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_2_io_to_pes_13_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_2_io_to_pes_14_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_2_io_to_pes_14_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_2_io_to_mem_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_2_io_to_mem_bits; // @[pe.scala 227:13]
  wire  PENetwork_3_io_to_pes_0_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_3_io_to_pes_0_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_3_io_to_pes_0_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_3_io_to_pes_0_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_3_io_to_pes_1_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_3_io_to_pes_1_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_3_io_to_pes_1_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_3_io_to_pes_1_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_3_io_to_pes_2_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_3_io_to_pes_2_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_3_io_to_pes_2_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_3_io_to_pes_2_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_3_io_to_pes_3_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_3_io_to_pes_3_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_3_io_to_pes_3_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_3_io_to_pes_3_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_3_io_to_pes_4_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_3_io_to_pes_4_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_3_io_to_pes_4_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_3_io_to_pes_4_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_3_io_to_pes_5_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_3_io_to_pes_5_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_3_io_to_pes_5_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_3_io_to_pes_5_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_3_io_to_pes_6_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_3_io_to_pes_6_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_3_io_to_pes_6_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_3_io_to_pes_6_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_3_io_to_pes_7_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_3_io_to_pes_7_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_3_io_to_pes_7_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_3_io_to_pes_7_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_3_io_to_pes_8_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_3_io_to_pes_8_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_3_io_to_pes_8_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_3_io_to_pes_8_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_3_io_to_pes_9_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_3_io_to_pes_9_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_3_io_to_pes_9_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_3_io_to_pes_9_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_3_io_to_pes_10_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_3_io_to_pes_10_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_3_io_to_pes_10_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_3_io_to_pes_10_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_3_io_to_pes_11_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_3_io_to_pes_11_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_3_io_to_pes_11_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_3_io_to_pes_11_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_3_io_to_pes_12_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_3_io_to_pes_12_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_3_io_to_pes_12_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_3_io_to_pes_12_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_3_io_to_pes_13_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_3_io_to_pes_13_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_3_io_to_pes_13_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_3_io_to_pes_13_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_3_io_to_pes_14_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_3_io_to_pes_14_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_3_io_to_mem_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_3_io_to_mem_bits; // @[pe.scala 227:13]
  wire  PENetwork_4_io_to_pes_0_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_4_io_to_pes_0_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_4_io_to_pes_0_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_4_io_to_pes_0_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_4_io_to_pes_1_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_4_io_to_pes_1_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_4_io_to_pes_1_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_4_io_to_pes_1_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_4_io_to_pes_2_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_4_io_to_pes_2_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_4_io_to_pes_2_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_4_io_to_pes_2_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_4_io_to_pes_3_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_4_io_to_pes_3_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_4_io_to_pes_3_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_4_io_to_pes_3_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_4_io_to_pes_4_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_4_io_to_pes_4_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_4_io_to_pes_4_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_4_io_to_pes_4_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_4_io_to_pes_5_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_4_io_to_pes_5_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_4_io_to_pes_5_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_4_io_to_pes_5_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_4_io_to_pes_6_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_4_io_to_pes_6_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_4_io_to_pes_6_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_4_io_to_pes_6_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_4_io_to_pes_7_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_4_io_to_pes_7_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_4_io_to_pes_7_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_4_io_to_pes_7_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_4_io_to_pes_8_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_4_io_to_pes_8_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_4_io_to_pes_8_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_4_io_to_pes_8_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_4_io_to_pes_9_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_4_io_to_pes_9_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_4_io_to_pes_9_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_4_io_to_pes_9_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_4_io_to_pes_10_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_4_io_to_pes_10_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_4_io_to_pes_10_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_4_io_to_pes_10_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_4_io_to_pes_11_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_4_io_to_pes_11_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_4_io_to_pes_11_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_4_io_to_pes_11_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_4_io_to_pes_12_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_4_io_to_pes_12_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_4_io_to_pes_12_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_4_io_to_pes_12_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_4_io_to_pes_13_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_4_io_to_pes_13_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_4_io_to_pes_13_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_4_io_to_pes_13_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_4_io_to_pes_14_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_4_io_to_pes_14_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_4_io_to_mem_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_4_io_to_mem_bits; // @[pe.scala 227:13]
  wire  PENetwork_5_io_to_pes_0_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_5_io_to_pes_0_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_5_io_to_pes_0_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_5_io_to_pes_0_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_5_io_to_pes_1_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_5_io_to_pes_1_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_5_io_to_pes_1_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_5_io_to_pes_1_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_5_io_to_pes_2_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_5_io_to_pes_2_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_5_io_to_pes_2_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_5_io_to_pes_2_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_5_io_to_pes_3_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_5_io_to_pes_3_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_5_io_to_pes_3_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_5_io_to_pes_3_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_5_io_to_pes_4_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_5_io_to_pes_4_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_5_io_to_pes_4_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_5_io_to_pes_4_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_5_io_to_pes_5_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_5_io_to_pes_5_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_5_io_to_pes_5_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_5_io_to_pes_5_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_5_io_to_pes_6_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_5_io_to_pes_6_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_5_io_to_pes_6_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_5_io_to_pes_6_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_5_io_to_pes_7_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_5_io_to_pes_7_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_5_io_to_pes_7_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_5_io_to_pes_7_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_5_io_to_pes_8_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_5_io_to_pes_8_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_5_io_to_pes_8_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_5_io_to_pes_8_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_5_io_to_pes_9_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_5_io_to_pes_9_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_5_io_to_pes_9_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_5_io_to_pes_9_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_5_io_to_pes_10_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_5_io_to_pes_10_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_5_io_to_pes_10_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_5_io_to_pes_10_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_5_io_to_pes_11_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_5_io_to_pes_11_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_5_io_to_pes_11_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_5_io_to_pes_11_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_5_io_to_pes_12_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_5_io_to_pes_12_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_5_io_to_pes_12_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_5_io_to_pes_12_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_5_io_to_pes_13_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_5_io_to_pes_13_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_5_io_to_pes_13_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_5_io_to_pes_13_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_5_io_to_pes_14_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_5_io_to_pes_14_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_5_io_to_mem_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_5_io_to_mem_bits; // @[pe.scala 227:13]
  wire  PENetwork_6_io_to_pes_0_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_6_io_to_pes_0_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_6_io_to_pes_0_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_6_io_to_pes_0_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_6_io_to_pes_1_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_6_io_to_pes_1_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_6_io_to_pes_1_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_6_io_to_pes_1_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_6_io_to_pes_2_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_6_io_to_pes_2_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_6_io_to_pes_2_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_6_io_to_pes_2_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_6_io_to_pes_3_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_6_io_to_pes_3_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_6_io_to_pes_3_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_6_io_to_pes_3_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_6_io_to_pes_4_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_6_io_to_pes_4_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_6_io_to_pes_4_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_6_io_to_pes_4_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_6_io_to_pes_5_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_6_io_to_pes_5_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_6_io_to_pes_5_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_6_io_to_pes_5_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_6_io_to_pes_6_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_6_io_to_pes_6_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_6_io_to_pes_6_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_6_io_to_pes_6_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_6_io_to_pes_7_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_6_io_to_pes_7_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_6_io_to_pes_7_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_6_io_to_pes_7_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_6_io_to_pes_8_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_6_io_to_pes_8_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_6_io_to_pes_8_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_6_io_to_pes_8_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_6_io_to_pes_9_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_6_io_to_pes_9_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_6_io_to_pes_9_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_6_io_to_pes_9_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_6_io_to_pes_10_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_6_io_to_pes_10_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_6_io_to_pes_10_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_6_io_to_pes_10_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_6_io_to_pes_11_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_6_io_to_pes_11_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_6_io_to_pes_11_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_6_io_to_pes_11_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_6_io_to_pes_12_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_6_io_to_pes_12_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_6_io_to_pes_12_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_6_io_to_pes_12_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_6_io_to_pes_13_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_6_io_to_pes_13_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_6_io_to_pes_13_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_6_io_to_pes_13_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_6_io_to_pes_14_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_6_io_to_pes_14_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_6_io_to_mem_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_6_io_to_mem_bits; // @[pe.scala 227:13]
  wire  PENetwork_7_io_to_pes_0_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_7_io_to_pes_0_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_7_io_to_pes_0_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_7_io_to_pes_0_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_7_io_to_pes_1_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_7_io_to_pes_1_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_7_io_to_pes_1_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_7_io_to_pes_1_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_7_io_to_pes_2_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_7_io_to_pes_2_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_7_io_to_pes_2_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_7_io_to_pes_2_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_7_io_to_pes_3_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_7_io_to_pes_3_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_7_io_to_pes_3_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_7_io_to_pes_3_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_7_io_to_pes_4_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_7_io_to_pes_4_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_7_io_to_pes_4_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_7_io_to_pes_4_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_7_io_to_pes_5_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_7_io_to_pes_5_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_7_io_to_pes_5_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_7_io_to_pes_5_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_7_io_to_pes_6_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_7_io_to_pes_6_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_7_io_to_pes_6_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_7_io_to_pes_6_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_7_io_to_pes_7_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_7_io_to_pes_7_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_7_io_to_pes_7_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_7_io_to_pes_7_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_7_io_to_pes_8_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_7_io_to_pes_8_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_7_io_to_pes_8_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_7_io_to_pes_8_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_7_io_to_pes_9_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_7_io_to_pes_9_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_7_io_to_pes_9_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_7_io_to_pes_9_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_7_io_to_pes_10_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_7_io_to_pes_10_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_7_io_to_pes_10_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_7_io_to_pes_10_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_7_io_to_pes_11_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_7_io_to_pes_11_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_7_io_to_pes_11_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_7_io_to_pes_11_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_7_io_to_pes_12_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_7_io_to_pes_12_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_7_io_to_pes_12_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_7_io_to_pes_12_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_7_io_to_pes_13_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_7_io_to_pes_13_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_7_io_to_pes_13_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_7_io_to_pes_13_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_7_io_to_pes_14_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_7_io_to_pes_14_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_7_io_to_mem_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_7_io_to_mem_bits; // @[pe.scala 227:13]
  wire  PENetwork_8_io_to_pes_0_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_8_io_to_pes_0_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_8_io_to_pes_0_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_8_io_to_pes_0_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_8_io_to_pes_1_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_8_io_to_pes_1_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_8_io_to_pes_1_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_8_io_to_pes_1_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_8_io_to_pes_2_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_8_io_to_pes_2_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_8_io_to_pes_2_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_8_io_to_pes_2_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_8_io_to_pes_3_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_8_io_to_pes_3_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_8_io_to_pes_3_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_8_io_to_pes_3_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_8_io_to_pes_4_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_8_io_to_pes_4_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_8_io_to_pes_4_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_8_io_to_pes_4_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_8_io_to_pes_5_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_8_io_to_pes_5_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_8_io_to_pes_5_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_8_io_to_pes_5_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_8_io_to_pes_6_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_8_io_to_pes_6_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_8_io_to_pes_6_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_8_io_to_pes_6_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_8_io_to_pes_7_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_8_io_to_pes_7_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_8_io_to_pes_7_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_8_io_to_pes_7_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_8_io_to_pes_8_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_8_io_to_pes_8_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_8_io_to_pes_8_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_8_io_to_pes_8_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_8_io_to_pes_9_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_8_io_to_pes_9_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_8_io_to_pes_9_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_8_io_to_pes_9_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_8_io_to_pes_10_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_8_io_to_pes_10_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_8_io_to_pes_10_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_8_io_to_pes_10_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_8_io_to_pes_11_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_8_io_to_pes_11_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_8_io_to_pes_11_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_8_io_to_pes_11_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_8_io_to_pes_12_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_8_io_to_pes_12_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_8_io_to_pes_12_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_8_io_to_pes_12_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_8_io_to_pes_13_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_8_io_to_pes_13_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_8_io_to_pes_13_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_8_io_to_pes_13_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_8_io_to_pes_14_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_8_io_to_pes_14_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_8_io_to_mem_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_8_io_to_mem_bits; // @[pe.scala 227:13]
  wire  PENetwork_9_io_to_pes_0_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_9_io_to_pes_0_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_9_io_to_pes_0_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_9_io_to_pes_0_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_9_io_to_pes_1_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_9_io_to_pes_1_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_9_io_to_pes_1_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_9_io_to_pes_1_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_9_io_to_pes_2_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_9_io_to_pes_2_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_9_io_to_pes_2_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_9_io_to_pes_2_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_9_io_to_pes_3_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_9_io_to_pes_3_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_9_io_to_pes_3_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_9_io_to_pes_3_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_9_io_to_pes_4_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_9_io_to_pes_4_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_9_io_to_pes_4_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_9_io_to_pes_4_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_9_io_to_pes_5_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_9_io_to_pes_5_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_9_io_to_pes_5_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_9_io_to_pes_5_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_9_io_to_pes_6_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_9_io_to_pes_6_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_9_io_to_pes_6_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_9_io_to_pes_6_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_9_io_to_pes_7_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_9_io_to_pes_7_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_9_io_to_pes_7_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_9_io_to_pes_7_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_9_io_to_pes_8_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_9_io_to_pes_8_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_9_io_to_pes_8_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_9_io_to_pes_8_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_9_io_to_pes_9_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_9_io_to_pes_9_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_9_io_to_pes_9_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_9_io_to_pes_9_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_9_io_to_pes_10_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_9_io_to_pes_10_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_9_io_to_pes_10_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_9_io_to_pes_10_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_9_io_to_pes_11_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_9_io_to_pes_11_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_9_io_to_pes_11_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_9_io_to_pes_11_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_9_io_to_pes_12_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_9_io_to_pes_12_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_9_io_to_pes_12_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_9_io_to_pes_12_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_9_io_to_pes_13_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_9_io_to_pes_13_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_9_io_to_pes_13_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_9_io_to_pes_13_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_9_io_to_pes_14_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_9_io_to_pes_14_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_9_io_to_mem_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_9_io_to_mem_bits; // @[pe.scala 227:13]
  wire  PENetwork_10_io_to_pes_0_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_10_io_to_pes_0_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_10_io_to_pes_0_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_10_io_to_pes_0_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_10_io_to_pes_1_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_10_io_to_pes_1_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_10_io_to_pes_1_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_10_io_to_pes_1_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_10_io_to_pes_2_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_10_io_to_pes_2_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_10_io_to_pes_2_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_10_io_to_pes_2_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_10_io_to_pes_3_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_10_io_to_pes_3_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_10_io_to_pes_3_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_10_io_to_pes_3_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_10_io_to_pes_4_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_10_io_to_pes_4_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_10_io_to_pes_4_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_10_io_to_pes_4_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_10_io_to_pes_5_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_10_io_to_pes_5_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_10_io_to_pes_5_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_10_io_to_pes_5_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_10_io_to_pes_6_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_10_io_to_pes_6_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_10_io_to_pes_6_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_10_io_to_pes_6_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_10_io_to_pes_7_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_10_io_to_pes_7_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_10_io_to_pes_7_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_10_io_to_pes_7_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_10_io_to_pes_8_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_10_io_to_pes_8_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_10_io_to_pes_8_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_10_io_to_pes_8_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_10_io_to_pes_9_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_10_io_to_pes_9_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_10_io_to_pes_9_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_10_io_to_pes_9_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_10_io_to_pes_10_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_10_io_to_pes_10_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_10_io_to_pes_10_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_10_io_to_pes_10_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_10_io_to_pes_11_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_10_io_to_pes_11_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_10_io_to_pes_11_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_10_io_to_pes_11_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_10_io_to_pes_12_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_10_io_to_pes_12_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_10_io_to_pes_12_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_10_io_to_pes_12_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_10_io_to_pes_13_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_10_io_to_pes_13_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_10_io_to_pes_13_out_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_10_io_to_pes_13_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_10_io_to_pes_14_in_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_10_io_to_pes_14_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_10_io_to_mem_valid; // @[pe.scala 227:13]
  wire [31:0] PENetwork_10_io_to_mem_bits; // @[pe.scala 227:13]
  wire  PENetwork_11_io_to_pes_0_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_11_io_to_pes_0_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_11_io_to_pes_0_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_11_io_to_pes_0_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_11_io_to_pes_1_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_11_io_to_pes_1_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_11_io_to_pes_1_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_11_io_to_pes_1_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_11_io_to_pes_2_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_11_io_to_pes_2_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_11_io_to_pes_2_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_11_io_to_pes_2_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_11_io_to_pes_3_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_11_io_to_pes_3_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_11_io_to_pes_3_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_11_io_to_pes_3_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_11_io_to_pes_4_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_11_io_to_pes_4_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_11_io_to_pes_4_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_11_io_to_pes_4_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_11_io_to_pes_5_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_11_io_to_pes_5_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_11_io_to_pes_5_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_11_io_to_pes_5_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_11_io_to_pes_6_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_11_io_to_pes_6_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_11_io_to_pes_6_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_11_io_to_pes_6_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_11_io_to_pes_7_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_11_io_to_pes_7_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_11_io_to_pes_7_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_11_io_to_pes_7_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_11_io_to_pes_8_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_11_io_to_pes_8_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_11_io_to_pes_8_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_11_io_to_pes_8_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_11_io_to_pes_9_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_11_io_to_pes_9_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_11_io_to_pes_9_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_11_io_to_pes_9_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_11_io_to_pes_10_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_11_io_to_pes_10_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_11_io_to_mem_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_11_io_to_mem_bits; // @[pe.scala 227:13]
  wire  PENetwork_12_io_to_pes_0_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_12_io_to_pes_0_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_12_io_to_pes_0_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_12_io_to_pes_0_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_12_io_to_pes_1_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_12_io_to_pes_1_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_12_io_to_pes_1_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_12_io_to_pes_1_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_12_io_to_pes_2_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_12_io_to_pes_2_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_12_io_to_pes_2_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_12_io_to_pes_2_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_12_io_to_pes_3_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_12_io_to_pes_3_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_12_io_to_pes_3_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_12_io_to_pes_3_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_12_io_to_pes_4_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_12_io_to_pes_4_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_12_io_to_pes_4_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_12_io_to_pes_4_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_12_io_to_pes_5_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_12_io_to_pes_5_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_12_io_to_pes_5_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_12_io_to_pes_5_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_12_io_to_pes_6_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_12_io_to_pes_6_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_12_io_to_pes_6_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_12_io_to_pes_6_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_12_io_to_pes_7_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_12_io_to_pes_7_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_12_io_to_pes_7_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_12_io_to_pes_7_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_12_io_to_pes_8_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_12_io_to_pes_8_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_12_io_to_pes_8_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_12_io_to_pes_8_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_12_io_to_pes_9_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_12_io_to_pes_9_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_12_io_to_pes_9_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_12_io_to_pes_9_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_12_io_to_pes_10_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_12_io_to_pes_10_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_12_io_to_mem_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_12_io_to_mem_bits; // @[pe.scala 227:13]
  wire  PENetwork_13_io_to_pes_0_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_13_io_to_pes_0_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_13_io_to_pes_0_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_13_io_to_pes_0_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_13_io_to_pes_1_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_13_io_to_pes_1_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_13_io_to_pes_1_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_13_io_to_pes_1_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_13_io_to_pes_2_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_13_io_to_pes_2_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_13_io_to_pes_2_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_13_io_to_pes_2_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_13_io_to_pes_3_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_13_io_to_pes_3_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_13_io_to_pes_3_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_13_io_to_pes_3_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_13_io_to_pes_4_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_13_io_to_pes_4_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_13_io_to_pes_4_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_13_io_to_pes_4_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_13_io_to_pes_5_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_13_io_to_pes_5_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_13_io_to_pes_5_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_13_io_to_pes_5_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_13_io_to_pes_6_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_13_io_to_pes_6_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_13_io_to_pes_6_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_13_io_to_pes_6_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_13_io_to_pes_7_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_13_io_to_pes_7_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_13_io_to_pes_7_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_13_io_to_pes_7_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_13_io_to_pes_8_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_13_io_to_pes_8_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_13_io_to_pes_8_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_13_io_to_pes_8_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_13_io_to_pes_9_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_13_io_to_pes_9_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_13_io_to_pes_9_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_13_io_to_pes_9_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_13_io_to_pes_10_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_13_io_to_pes_10_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_13_io_to_mem_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_13_io_to_mem_bits; // @[pe.scala 227:13]
  wire  PENetwork_14_io_to_pes_0_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_14_io_to_pes_0_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_14_io_to_pes_0_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_14_io_to_pes_0_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_14_io_to_pes_1_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_14_io_to_pes_1_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_14_io_to_pes_1_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_14_io_to_pes_1_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_14_io_to_pes_2_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_14_io_to_pes_2_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_14_io_to_pes_2_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_14_io_to_pes_2_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_14_io_to_pes_3_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_14_io_to_pes_3_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_14_io_to_pes_3_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_14_io_to_pes_3_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_14_io_to_pes_4_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_14_io_to_pes_4_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_14_io_to_pes_4_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_14_io_to_pes_4_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_14_io_to_pes_5_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_14_io_to_pes_5_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_14_io_to_pes_5_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_14_io_to_pes_5_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_14_io_to_pes_6_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_14_io_to_pes_6_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_14_io_to_pes_6_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_14_io_to_pes_6_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_14_io_to_pes_7_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_14_io_to_pes_7_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_14_io_to_pes_7_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_14_io_to_pes_7_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_14_io_to_pes_8_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_14_io_to_pes_8_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_14_io_to_pes_8_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_14_io_to_pes_8_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_14_io_to_pes_9_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_14_io_to_pes_9_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_14_io_to_pes_9_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_14_io_to_pes_9_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_14_io_to_pes_10_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_14_io_to_pes_10_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_14_io_to_mem_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_14_io_to_mem_bits; // @[pe.scala 227:13]
  wire  PENetwork_15_io_to_pes_0_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_15_io_to_pes_0_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_15_io_to_pes_0_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_15_io_to_pes_0_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_15_io_to_pes_1_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_15_io_to_pes_1_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_15_io_to_pes_1_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_15_io_to_pes_1_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_15_io_to_pes_2_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_15_io_to_pes_2_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_15_io_to_pes_2_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_15_io_to_pes_2_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_15_io_to_pes_3_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_15_io_to_pes_3_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_15_io_to_pes_3_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_15_io_to_pes_3_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_15_io_to_pes_4_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_15_io_to_pes_4_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_15_io_to_pes_4_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_15_io_to_pes_4_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_15_io_to_pes_5_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_15_io_to_pes_5_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_15_io_to_pes_5_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_15_io_to_pes_5_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_15_io_to_pes_6_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_15_io_to_pes_6_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_15_io_to_pes_6_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_15_io_to_pes_6_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_15_io_to_pes_7_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_15_io_to_pes_7_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_15_io_to_pes_7_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_15_io_to_pes_7_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_15_io_to_pes_8_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_15_io_to_pes_8_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_15_io_to_pes_8_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_15_io_to_pes_8_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_15_io_to_pes_9_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_15_io_to_pes_9_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_15_io_to_pes_9_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_15_io_to_pes_9_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_15_io_to_pes_10_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_15_io_to_pes_10_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_15_io_to_mem_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_15_io_to_mem_bits; // @[pe.scala 227:13]
  wire  PENetwork_16_io_to_pes_0_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_16_io_to_pes_0_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_16_io_to_pes_0_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_16_io_to_pes_0_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_16_io_to_pes_1_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_16_io_to_pes_1_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_16_io_to_pes_1_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_16_io_to_pes_1_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_16_io_to_pes_2_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_16_io_to_pes_2_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_16_io_to_pes_2_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_16_io_to_pes_2_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_16_io_to_pes_3_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_16_io_to_pes_3_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_16_io_to_pes_3_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_16_io_to_pes_3_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_16_io_to_pes_4_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_16_io_to_pes_4_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_16_io_to_pes_4_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_16_io_to_pes_4_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_16_io_to_pes_5_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_16_io_to_pes_5_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_16_io_to_pes_5_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_16_io_to_pes_5_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_16_io_to_pes_6_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_16_io_to_pes_6_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_16_io_to_pes_6_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_16_io_to_pes_6_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_16_io_to_pes_7_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_16_io_to_pes_7_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_16_io_to_pes_7_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_16_io_to_pes_7_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_16_io_to_pes_8_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_16_io_to_pes_8_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_16_io_to_pes_8_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_16_io_to_pes_8_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_16_io_to_pes_9_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_16_io_to_pes_9_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_16_io_to_pes_9_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_16_io_to_pes_9_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_16_io_to_pes_10_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_16_io_to_pes_10_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_16_io_to_mem_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_16_io_to_mem_bits; // @[pe.scala 227:13]
  wire  PENetwork_17_io_to_pes_0_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_17_io_to_pes_0_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_17_io_to_pes_0_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_17_io_to_pes_0_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_17_io_to_pes_1_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_17_io_to_pes_1_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_17_io_to_pes_1_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_17_io_to_pes_1_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_17_io_to_pes_2_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_17_io_to_pes_2_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_17_io_to_pes_2_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_17_io_to_pes_2_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_17_io_to_pes_3_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_17_io_to_pes_3_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_17_io_to_pes_3_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_17_io_to_pes_3_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_17_io_to_pes_4_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_17_io_to_pes_4_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_17_io_to_pes_4_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_17_io_to_pes_4_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_17_io_to_pes_5_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_17_io_to_pes_5_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_17_io_to_pes_5_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_17_io_to_pes_5_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_17_io_to_pes_6_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_17_io_to_pes_6_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_17_io_to_pes_6_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_17_io_to_pes_6_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_17_io_to_pes_7_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_17_io_to_pes_7_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_17_io_to_pes_7_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_17_io_to_pes_7_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_17_io_to_pes_8_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_17_io_to_pes_8_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_17_io_to_pes_8_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_17_io_to_pes_8_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_17_io_to_pes_9_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_17_io_to_pes_9_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_17_io_to_pes_9_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_17_io_to_pes_9_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_17_io_to_pes_10_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_17_io_to_pes_10_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_17_io_to_mem_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_17_io_to_mem_bits; // @[pe.scala 227:13]
  wire  PENetwork_18_io_to_pes_0_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_18_io_to_pes_0_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_18_io_to_pes_0_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_18_io_to_pes_0_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_18_io_to_pes_1_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_18_io_to_pes_1_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_18_io_to_pes_1_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_18_io_to_pes_1_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_18_io_to_pes_2_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_18_io_to_pes_2_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_18_io_to_pes_2_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_18_io_to_pes_2_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_18_io_to_pes_3_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_18_io_to_pes_3_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_18_io_to_pes_3_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_18_io_to_pes_3_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_18_io_to_pes_4_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_18_io_to_pes_4_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_18_io_to_pes_4_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_18_io_to_pes_4_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_18_io_to_pes_5_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_18_io_to_pes_5_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_18_io_to_pes_5_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_18_io_to_pes_5_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_18_io_to_pes_6_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_18_io_to_pes_6_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_18_io_to_pes_6_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_18_io_to_pes_6_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_18_io_to_pes_7_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_18_io_to_pes_7_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_18_io_to_pes_7_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_18_io_to_pes_7_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_18_io_to_pes_8_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_18_io_to_pes_8_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_18_io_to_pes_8_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_18_io_to_pes_8_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_18_io_to_pes_9_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_18_io_to_pes_9_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_18_io_to_pes_9_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_18_io_to_pes_9_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_18_io_to_pes_10_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_18_io_to_pes_10_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_18_io_to_mem_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_18_io_to_mem_bits; // @[pe.scala 227:13]
  wire  PENetwork_19_io_to_pes_0_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_19_io_to_pes_0_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_19_io_to_pes_0_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_19_io_to_pes_0_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_19_io_to_pes_1_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_19_io_to_pes_1_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_19_io_to_pes_1_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_19_io_to_pes_1_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_19_io_to_pes_2_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_19_io_to_pes_2_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_19_io_to_pes_2_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_19_io_to_pes_2_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_19_io_to_pes_3_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_19_io_to_pes_3_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_19_io_to_pes_3_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_19_io_to_pes_3_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_19_io_to_pes_4_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_19_io_to_pes_4_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_19_io_to_pes_4_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_19_io_to_pes_4_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_19_io_to_pes_5_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_19_io_to_pes_5_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_19_io_to_pes_5_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_19_io_to_pes_5_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_19_io_to_pes_6_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_19_io_to_pes_6_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_19_io_to_pes_6_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_19_io_to_pes_6_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_19_io_to_pes_7_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_19_io_to_pes_7_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_19_io_to_pes_7_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_19_io_to_pes_7_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_19_io_to_pes_8_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_19_io_to_pes_8_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_19_io_to_pes_8_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_19_io_to_pes_8_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_19_io_to_pes_9_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_19_io_to_pes_9_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_19_io_to_pes_9_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_19_io_to_pes_9_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_19_io_to_pes_10_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_19_io_to_pes_10_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_19_io_to_mem_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_19_io_to_mem_bits; // @[pe.scala 227:13]
  wire  PENetwork_20_io_to_pes_0_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_20_io_to_pes_0_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_20_io_to_pes_0_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_20_io_to_pes_0_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_20_io_to_pes_1_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_20_io_to_pes_1_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_20_io_to_pes_1_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_20_io_to_pes_1_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_20_io_to_pes_2_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_20_io_to_pes_2_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_20_io_to_pes_2_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_20_io_to_pes_2_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_20_io_to_pes_3_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_20_io_to_pes_3_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_20_io_to_pes_3_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_20_io_to_pes_3_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_20_io_to_pes_4_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_20_io_to_pes_4_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_20_io_to_pes_4_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_20_io_to_pes_4_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_20_io_to_pes_5_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_20_io_to_pes_5_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_20_io_to_pes_5_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_20_io_to_pes_5_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_20_io_to_pes_6_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_20_io_to_pes_6_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_20_io_to_pes_6_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_20_io_to_pes_6_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_20_io_to_pes_7_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_20_io_to_pes_7_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_20_io_to_pes_7_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_20_io_to_pes_7_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_20_io_to_pes_8_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_20_io_to_pes_8_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_20_io_to_pes_8_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_20_io_to_pes_8_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_20_io_to_pes_9_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_20_io_to_pes_9_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_20_io_to_pes_9_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_20_io_to_pes_9_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_20_io_to_pes_10_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_20_io_to_pes_10_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_20_io_to_mem_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_20_io_to_mem_bits; // @[pe.scala 227:13]
  wire  PENetwork_21_io_to_pes_0_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_21_io_to_pes_0_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_21_io_to_pes_0_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_21_io_to_pes_0_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_21_io_to_pes_1_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_21_io_to_pes_1_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_21_io_to_pes_1_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_21_io_to_pes_1_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_21_io_to_pes_2_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_21_io_to_pes_2_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_21_io_to_pes_2_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_21_io_to_pes_2_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_21_io_to_pes_3_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_21_io_to_pes_3_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_21_io_to_pes_3_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_21_io_to_pes_3_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_21_io_to_pes_4_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_21_io_to_pes_4_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_21_io_to_pes_4_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_21_io_to_pes_4_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_21_io_to_pes_5_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_21_io_to_pes_5_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_21_io_to_pes_5_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_21_io_to_pes_5_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_21_io_to_pes_6_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_21_io_to_pes_6_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_21_io_to_pes_6_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_21_io_to_pes_6_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_21_io_to_pes_7_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_21_io_to_pes_7_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_21_io_to_pes_7_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_21_io_to_pes_7_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_21_io_to_pes_8_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_21_io_to_pes_8_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_21_io_to_pes_8_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_21_io_to_pes_8_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_21_io_to_pes_9_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_21_io_to_pes_9_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_21_io_to_pes_9_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_21_io_to_pes_9_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_21_io_to_pes_10_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_21_io_to_pes_10_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_21_io_to_mem_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_21_io_to_mem_bits; // @[pe.scala 227:13]
  wire  PENetwork_22_io_to_pes_0_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_22_io_to_pes_0_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_22_io_to_pes_0_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_22_io_to_pes_0_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_22_io_to_pes_1_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_22_io_to_pes_1_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_22_io_to_pes_1_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_22_io_to_pes_1_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_22_io_to_pes_2_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_22_io_to_pes_2_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_22_io_to_pes_2_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_22_io_to_pes_2_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_22_io_to_pes_3_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_22_io_to_pes_3_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_22_io_to_pes_3_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_22_io_to_pes_3_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_22_io_to_pes_4_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_22_io_to_pes_4_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_22_io_to_pes_4_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_22_io_to_pes_4_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_22_io_to_pes_5_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_22_io_to_pes_5_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_22_io_to_pes_5_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_22_io_to_pes_5_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_22_io_to_pes_6_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_22_io_to_pes_6_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_22_io_to_pes_6_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_22_io_to_pes_6_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_22_io_to_pes_7_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_22_io_to_pes_7_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_22_io_to_pes_7_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_22_io_to_pes_7_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_22_io_to_pes_8_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_22_io_to_pes_8_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_22_io_to_pes_8_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_22_io_to_pes_8_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_22_io_to_pes_9_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_22_io_to_pes_9_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_22_io_to_pes_9_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_22_io_to_pes_9_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_22_io_to_pes_10_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_22_io_to_pes_10_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_22_io_to_mem_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_22_io_to_mem_bits; // @[pe.scala 227:13]
  wire  PENetwork_23_io_to_pes_0_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_23_io_to_pes_0_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_23_io_to_pes_0_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_23_io_to_pes_0_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_23_io_to_pes_1_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_23_io_to_pes_1_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_23_io_to_pes_1_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_23_io_to_pes_1_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_23_io_to_pes_2_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_23_io_to_pes_2_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_23_io_to_pes_2_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_23_io_to_pes_2_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_23_io_to_pes_3_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_23_io_to_pes_3_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_23_io_to_pes_3_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_23_io_to_pes_3_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_23_io_to_pes_4_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_23_io_to_pes_4_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_23_io_to_pes_4_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_23_io_to_pes_4_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_23_io_to_pes_5_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_23_io_to_pes_5_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_23_io_to_pes_5_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_23_io_to_pes_5_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_23_io_to_pes_6_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_23_io_to_pes_6_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_23_io_to_pes_6_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_23_io_to_pes_6_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_23_io_to_pes_7_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_23_io_to_pes_7_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_23_io_to_pes_7_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_23_io_to_pes_7_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_23_io_to_pes_8_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_23_io_to_pes_8_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_23_io_to_pes_8_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_23_io_to_pes_8_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_23_io_to_pes_9_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_23_io_to_pes_9_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_23_io_to_pes_9_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_23_io_to_pes_9_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_23_io_to_pes_10_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_23_io_to_pes_10_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_23_io_to_mem_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_23_io_to_mem_bits; // @[pe.scala 227:13]
  wire  PENetwork_24_io_to_pes_0_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_24_io_to_pes_0_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_24_io_to_pes_0_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_24_io_to_pes_0_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_24_io_to_pes_1_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_24_io_to_pes_1_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_24_io_to_pes_1_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_24_io_to_pes_1_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_24_io_to_pes_2_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_24_io_to_pes_2_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_24_io_to_pes_2_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_24_io_to_pes_2_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_24_io_to_pes_3_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_24_io_to_pes_3_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_24_io_to_pes_3_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_24_io_to_pes_3_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_24_io_to_pes_4_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_24_io_to_pes_4_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_24_io_to_pes_4_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_24_io_to_pes_4_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_24_io_to_pes_5_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_24_io_to_pes_5_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_24_io_to_pes_5_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_24_io_to_pes_5_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_24_io_to_pes_6_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_24_io_to_pes_6_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_24_io_to_pes_6_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_24_io_to_pes_6_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_24_io_to_pes_7_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_24_io_to_pes_7_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_24_io_to_pes_7_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_24_io_to_pes_7_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_24_io_to_pes_8_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_24_io_to_pes_8_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_24_io_to_pes_8_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_24_io_to_pes_8_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_24_io_to_pes_9_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_24_io_to_pes_9_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_24_io_to_pes_9_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_24_io_to_pes_9_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_24_io_to_pes_10_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_24_io_to_pes_10_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_24_io_to_mem_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_24_io_to_mem_bits; // @[pe.scala 227:13]
  wire  PENetwork_25_io_to_pes_0_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_25_io_to_pes_0_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_25_io_to_pes_0_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_25_io_to_pes_0_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_25_io_to_pes_1_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_25_io_to_pes_1_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_25_io_to_pes_1_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_25_io_to_pes_1_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_25_io_to_pes_2_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_25_io_to_pes_2_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_25_io_to_pes_2_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_25_io_to_pes_2_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_25_io_to_pes_3_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_25_io_to_pes_3_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_25_io_to_pes_3_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_25_io_to_pes_3_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_25_io_to_pes_4_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_25_io_to_pes_4_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_25_io_to_pes_4_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_25_io_to_pes_4_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_25_io_to_pes_5_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_25_io_to_pes_5_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_25_io_to_pes_5_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_25_io_to_pes_5_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_25_io_to_pes_6_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_25_io_to_pes_6_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_25_io_to_pes_6_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_25_io_to_pes_6_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_25_io_to_pes_7_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_25_io_to_pes_7_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_25_io_to_pes_7_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_25_io_to_pes_7_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_25_io_to_pes_8_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_25_io_to_pes_8_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_25_io_to_pes_8_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_25_io_to_pes_8_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_25_io_to_pes_9_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_25_io_to_pes_9_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_25_io_to_pes_9_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_25_io_to_pes_9_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_25_io_to_pes_10_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_25_io_to_pes_10_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_25_io_to_mem_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_25_io_to_mem_bits; // @[pe.scala 227:13]
  wire  PENetwork_26_clock; // @[pe.scala 227:13]
  wire  PENetwork_26_io_to_pes_0_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_26_io_to_pes_0_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_26_io_to_pes_0_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_26_io_to_pes_0_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_26_io_to_pes_1_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_26_io_to_pes_1_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_26_io_to_pes_1_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_26_io_to_pes_1_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_26_io_to_pes_1_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_26_io_to_pes_1_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_26_io_to_pes_1_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_26_io_to_pes_2_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_26_io_to_pes_2_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_26_io_to_pes_2_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_26_io_to_pes_2_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_26_io_to_pes_2_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_26_io_to_pes_2_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_26_io_to_pes_2_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_26_io_to_pes_3_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_26_io_to_pes_3_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_26_io_to_pes_3_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_26_io_to_pes_3_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_26_io_to_pes_3_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_26_io_to_pes_3_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_26_io_to_pes_3_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_26_io_to_pes_4_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_26_io_to_pes_4_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_26_io_to_pes_4_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_26_io_to_pes_4_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_26_io_to_pes_4_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_26_io_to_pes_4_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_26_io_to_pes_4_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_26_io_to_pes_5_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_26_io_to_pes_5_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_26_io_to_pes_5_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_26_io_to_pes_5_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_26_io_to_pes_5_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_26_io_to_pes_5_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_26_io_to_pes_5_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_26_io_to_pes_6_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_26_io_to_pes_6_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_26_io_to_pes_6_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_26_io_to_pes_6_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_26_io_to_pes_6_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_26_io_to_pes_6_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_26_io_to_pes_6_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_26_io_to_pes_7_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_26_io_to_pes_7_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_26_io_to_pes_7_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_26_io_to_pes_7_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_26_io_to_pes_7_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_26_io_to_pes_7_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_26_io_to_pes_7_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_26_io_to_pes_8_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_26_io_to_pes_8_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_26_io_to_pes_8_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_26_io_to_pes_8_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_26_io_to_pes_8_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_26_io_to_pes_8_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_26_io_to_pes_8_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_26_io_to_pes_9_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_26_io_to_pes_9_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_26_io_to_pes_9_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_26_io_to_pes_9_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_26_io_to_pes_9_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_26_io_to_pes_9_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_26_io_to_pes_9_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_26_io_to_pes_10_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_26_io_to_pes_10_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_26_io_to_pes_10_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_26_io_to_pes_10_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_26_io_to_pes_10_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_26_io_to_pes_10_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_26_io_to_mem_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_26_io_to_mem_bits; // @[pe.scala 227:13]
  wire  PENetwork_26_io_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_27_clock; // @[pe.scala 227:13]
  wire  PENetwork_27_io_to_pes_0_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_27_io_to_pes_0_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_27_io_to_pes_0_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_27_io_to_pes_0_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_27_io_to_pes_1_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_27_io_to_pes_1_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_27_io_to_pes_1_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_27_io_to_pes_1_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_27_io_to_pes_1_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_27_io_to_pes_1_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_27_io_to_pes_1_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_27_io_to_pes_2_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_27_io_to_pes_2_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_27_io_to_pes_2_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_27_io_to_pes_2_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_27_io_to_pes_2_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_27_io_to_pes_2_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_27_io_to_pes_2_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_27_io_to_pes_3_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_27_io_to_pes_3_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_27_io_to_pes_3_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_27_io_to_pes_3_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_27_io_to_pes_3_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_27_io_to_pes_3_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_27_io_to_pes_3_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_27_io_to_pes_4_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_27_io_to_pes_4_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_27_io_to_pes_4_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_27_io_to_pes_4_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_27_io_to_pes_4_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_27_io_to_pes_4_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_27_io_to_pes_4_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_27_io_to_pes_5_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_27_io_to_pes_5_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_27_io_to_pes_5_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_27_io_to_pes_5_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_27_io_to_pes_5_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_27_io_to_pes_5_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_27_io_to_pes_5_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_27_io_to_pes_6_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_27_io_to_pes_6_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_27_io_to_pes_6_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_27_io_to_pes_6_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_27_io_to_pes_6_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_27_io_to_pes_6_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_27_io_to_pes_6_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_27_io_to_pes_7_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_27_io_to_pes_7_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_27_io_to_pes_7_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_27_io_to_pes_7_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_27_io_to_pes_7_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_27_io_to_pes_7_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_27_io_to_pes_7_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_27_io_to_pes_8_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_27_io_to_pes_8_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_27_io_to_pes_8_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_27_io_to_pes_8_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_27_io_to_pes_8_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_27_io_to_pes_8_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_27_io_to_pes_8_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_27_io_to_pes_9_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_27_io_to_pes_9_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_27_io_to_pes_9_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_27_io_to_pes_9_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_27_io_to_pes_9_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_27_io_to_pes_9_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_27_io_to_pes_9_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_27_io_to_pes_10_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_27_io_to_pes_10_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_27_io_to_pes_10_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_27_io_to_pes_10_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_27_io_to_pes_10_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_27_io_to_pes_10_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_27_io_to_mem_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_27_io_to_mem_bits; // @[pe.scala 227:13]
  wire  PENetwork_27_io_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_28_clock; // @[pe.scala 227:13]
  wire  PENetwork_28_io_to_pes_0_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_28_io_to_pes_0_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_28_io_to_pes_0_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_28_io_to_pes_0_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_28_io_to_pes_1_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_28_io_to_pes_1_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_28_io_to_pes_1_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_28_io_to_pes_1_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_28_io_to_pes_1_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_28_io_to_pes_1_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_28_io_to_pes_1_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_28_io_to_pes_2_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_28_io_to_pes_2_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_28_io_to_pes_2_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_28_io_to_pes_2_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_28_io_to_pes_2_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_28_io_to_pes_2_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_28_io_to_pes_2_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_28_io_to_pes_3_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_28_io_to_pes_3_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_28_io_to_pes_3_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_28_io_to_pes_3_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_28_io_to_pes_3_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_28_io_to_pes_3_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_28_io_to_pes_3_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_28_io_to_pes_4_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_28_io_to_pes_4_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_28_io_to_pes_4_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_28_io_to_pes_4_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_28_io_to_pes_4_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_28_io_to_pes_4_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_28_io_to_pes_4_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_28_io_to_pes_5_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_28_io_to_pes_5_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_28_io_to_pes_5_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_28_io_to_pes_5_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_28_io_to_pes_5_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_28_io_to_pes_5_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_28_io_to_pes_5_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_28_io_to_pes_6_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_28_io_to_pes_6_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_28_io_to_pes_6_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_28_io_to_pes_6_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_28_io_to_pes_6_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_28_io_to_pes_6_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_28_io_to_pes_6_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_28_io_to_pes_7_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_28_io_to_pes_7_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_28_io_to_pes_7_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_28_io_to_pes_7_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_28_io_to_pes_7_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_28_io_to_pes_7_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_28_io_to_pes_7_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_28_io_to_pes_8_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_28_io_to_pes_8_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_28_io_to_pes_8_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_28_io_to_pes_8_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_28_io_to_pes_8_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_28_io_to_pes_8_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_28_io_to_pes_8_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_28_io_to_pes_9_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_28_io_to_pes_9_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_28_io_to_pes_9_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_28_io_to_pes_9_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_28_io_to_pes_9_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_28_io_to_pes_9_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_28_io_to_pes_9_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_28_io_to_pes_10_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_28_io_to_pes_10_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_28_io_to_pes_10_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_28_io_to_pes_10_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_28_io_to_pes_10_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_28_io_to_pes_10_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_28_io_to_mem_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_28_io_to_mem_bits; // @[pe.scala 227:13]
  wire  PENetwork_28_io_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_29_clock; // @[pe.scala 227:13]
  wire  PENetwork_29_io_to_pes_0_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_29_io_to_pes_0_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_29_io_to_pes_0_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_29_io_to_pes_0_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_29_io_to_pes_1_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_29_io_to_pes_1_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_29_io_to_pes_1_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_29_io_to_pes_1_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_29_io_to_pes_1_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_29_io_to_pes_1_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_29_io_to_pes_1_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_29_io_to_pes_2_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_29_io_to_pes_2_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_29_io_to_pes_2_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_29_io_to_pes_2_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_29_io_to_pes_2_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_29_io_to_pes_2_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_29_io_to_pes_2_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_29_io_to_pes_3_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_29_io_to_pes_3_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_29_io_to_pes_3_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_29_io_to_pes_3_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_29_io_to_pes_3_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_29_io_to_pes_3_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_29_io_to_pes_3_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_29_io_to_pes_4_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_29_io_to_pes_4_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_29_io_to_pes_4_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_29_io_to_pes_4_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_29_io_to_pes_4_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_29_io_to_pes_4_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_29_io_to_pes_4_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_29_io_to_pes_5_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_29_io_to_pes_5_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_29_io_to_pes_5_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_29_io_to_pes_5_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_29_io_to_pes_5_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_29_io_to_pes_5_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_29_io_to_pes_5_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_29_io_to_pes_6_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_29_io_to_pes_6_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_29_io_to_pes_6_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_29_io_to_pes_6_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_29_io_to_pes_6_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_29_io_to_pes_6_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_29_io_to_pes_6_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_29_io_to_pes_7_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_29_io_to_pes_7_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_29_io_to_pes_7_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_29_io_to_pes_7_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_29_io_to_pes_7_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_29_io_to_pes_7_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_29_io_to_pes_7_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_29_io_to_pes_8_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_29_io_to_pes_8_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_29_io_to_pes_8_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_29_io_to_pes_8_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_29_io_to_pes_8_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_29_io_to_pes_8_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_29_io_to_pes_8_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_29_io_to_pes_9_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_29_io_to_pes_9_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_29_io_to_pes_9_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_29_io_to_pes_9_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_29_io_to_pes_9_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_29_io_to_pes_9_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_29_io_to_pes_9_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_29_io_to_pes_10_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_29_io_to_pes_10_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_29_io_to_pes_10_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_29_io_to_pes_10_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_29_io_to_pes_10_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_29_io_to_pes_10_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_29_io_to_mem_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_29_io_to_mem_bits; // @[pe.scala 227:13]
  wire  PENetwork_29_io_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_30_clock; // @[pe.scala 227:13]
  wire  PENetwork_30_io_to_pes_0_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_30_io_to_pes_0_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_30_io_to_pes_0_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_30_io_to_pes_0_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_30_io_to_pes_1_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_30_io_to_pes_1_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_30_io_to_pes_1_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_30_io_to_pes_1_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_30_io_to_pes_1_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_30_io_to_pes_1_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_30_io_to_pes_1_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_30_io_to_pes_2_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_30_io_to_pes_2_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_30_io_to_pes_2_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_30_io_to_pes_2_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_30_io_to_pes_2_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_30_io_to_pes_2_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_30_io_to_pes_2_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_30_io_to_pes_3_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_30_io_to_pes_3_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_30_io_to_pes_3_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_30_io_to_pes_3_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_30_io_to_pes_3_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_30_io_to_pes_3_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_30_io_to_pes_3_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_30_io_to_pes_4_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_30_io_to_pes_4_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_30_io_to_pes_4_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_30_io_to_pes_4_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_30_io_to_pes_4_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_30_io_to_pes_4_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_30_io_to_pes_4_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_30_io_to_pes_5_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_30_io_to_pes_5_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_30_io_to_pes_5_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_30_io_to_pes_5_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_30_io_to_pes_5_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_30_io_to_pes_5_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_30_io_to_pes_5_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_30_io_to_pes_6_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_30_io_to_pes_6_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_30_io_to_pes_6_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_30_io_to_pes_6_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_30_io_to_pes_6_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_30_io_to_pes_6_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_30_io_to_pes_6_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_30_io_to_pes_7_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_30_io_to_pes_7_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_30_io_to_pes_7_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_30_io_to_pes_7_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_30_io_to_pes_7_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_30_io_to_pes_7_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_30_io_to_pes_7_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_30_io_to_pes_8_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_30_io_to_pes_8_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_30_io_to_pes_8_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_30_io_to_pes_8_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_30_io_to_pes_8_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_30_io_to_pes_8_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_30_io_to_pes_8_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_30_io_to_pes_9_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_30_io_to_pes_9_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_30_io_to_pes_9_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_30_io_to_pes_9_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_30_io_to_pes_9_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_30_io_to_pes_9_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_30_io_to_pes_9_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_30_io_to_pes_10_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_30_io_to_pes_10_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_30_io_to_pes_10_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_30_io_to_pes_10_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_30_io_to_pes_10_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_30_io_to_pes_10_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_30_io_to_mem_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_30_io_to_mem_bits; // @[pe.scala 227:13]
  wire  PENetwork_30_io_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_31_clock; // @[pe.scala 227:13]
  wire  PENetwork_31_io_to_pes_0_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_31_io_to_pes_0_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_31_io_to_pes_0_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_31_io_to_pes_0_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_31_io_to_pes_1_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_31_io_to_pes_1_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_31_io_to_pes_1_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_31_io_to_pes_1_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_31_io_to_pes_1_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_31_io_to_pes_1_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_31_io_to_pes_1_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_31_io_to_pes_2_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_31_io_to_pes_2_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_31_io_to_pes_2_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_31_io_to_pes_2_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_31_io_to_pes_2_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_31_io_to_pes_2_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_31_io_to_pes_2_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_31_io_to_pes_3_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_31_io_to_pes_3_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_31_io_to_pes_3_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_31_io_to_pes_3_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_31_io_to_pes_3_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_31_io_to_pes_3_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_31_io_to_pes_3_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_31_io_to_pes_4_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_31_io_to_pes_4_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_31_io_to_pes_4_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_31_io_to_pes_4_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_31_io_to_pes_4_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_31_io_to_pes_4_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_31_io_to_pes_4_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_31_io_to_pes_5_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_31_io_to_pes_5_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_31_io_to_pes_5_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_31_io_to_pes_5_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_31_io_to_pes_5_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_31_io_to_pes_5_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_31_io_to_pes_5_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_31_io_to_pes_6_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_31_io_to_pes_6_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_31_io_to_pes_6_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_31_io_to_pes_6_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_31_io_to_pes_6_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_31_io_to_pes_6_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_31_io_to_pes_6_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_31_io_to_pes_7_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_31_io_to_pes_7_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_31_io_to_pes_7_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_31_io_to_pes_7_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_31_io_to_pes_7_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_31_io_to_pes_7_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_31_io_to_pes_7_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_31_io_to_pes_8_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_31_io_to_pes_8_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_31_io_to_pes_8_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_31_io_to_pes_8_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_31_io_to_pes_8_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_31_io_to_pes_8_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_31_io_to_pes_8_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_31_io_to_pes_9_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_31_io_to_pes_9_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_31_io_to_pes_9_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_31_io_to_pes_9_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_31_io_to_pes_9_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_31_io_to_pes_9_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_31_io_to_pes_9_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_31_io_to_pes_10_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_31_io_to_pes_10_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_31_io_to_pes_10_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_31_io_to_pes_10_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_31_io_to_pes_10_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_31_io_to_pes_10_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_31_io_to_mem_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_31_io_to_mem_bits; // @[pe.scala 227:13]
  wire  PENetwork_31_io_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_32_clock; // @[pe.scala 227:13]
  wire  PENetwork_32_io_to_pes_0_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_32_io_to_pes_0_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_32_io_to_pes_0_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_32_io_to_pes_0_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_32_io_to_pes_1_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_32_io_to_pes_1_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_32_io_to_pes_1_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_32_io_to_pes_1_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_32_io_to_pes_1_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_32_io_to_pes_1_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_32_io_to_pes_1_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_32_io_to_pes_2_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_32_io_to_pes_2_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_32_io_to_pes_2_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_32_io_to_pes_2_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_32_io_to_pes_2_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_32_io_to_pes_2_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_32_io_to_pes_2_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_32_io_to_pes_3_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_32_io_to_pes_3_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_32_io_to_pes_3_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_32_io_to_pes_3_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_32_io_to_pes_3_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_32_io_to_pes_3_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_32_io_to_pes_3_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_32_io_to_pes_4_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_32_io_to_pes_4_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_32_io_to_pes_4_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_32_io_to_pes_4_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_32_io_to_pes_4_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_32_io_to_pes_4_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_32_io_to_pes_4_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_32_io_to_pes_5_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_32_io_to_pes_5_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_32_io_to_pes_5_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_32_io_to_pes_5_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_32_io_to_pes_5_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_32_io_to_pes_5_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_32_io_to_pes_5_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_32_io_to_pes_6_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_32_io_to_pes_6_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_32_io_to_pes_6_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_32_io_to_pes_6_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_32_io_to_pes_6_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_32_io_to_pes_6_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_32_io_to_pes_6_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_32_io_to_pes_7_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_32_io_to_pes_7_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_32_io_to_pes_7_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_32_io_to_pes_7_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_32_io_to_pes_7_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_32_io_to_pes_7_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_32_io_to_pes_7_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_32_io_to_pes_8_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_32_io_to_pes_8_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_32_io_to_pes_8_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_32_io_to_pes_8_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_32_io_to_pes_8_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_32_io_to_pes_8_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_32_io_to_pes_8_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_32_io_to_pes_9_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_32_io_to_pes_9_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_32_io_to_pes_9_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_32_io_to_pes_9_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_32_io_to_pes_9_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_32_io_to_pes_9_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_32_io_to_pes_9_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_32_io_to_pes_10_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_32_io_to_pes_10_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_32_io_to_pes_10_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_32_io_to_pes_10_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_32_io_to_pes_10_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_32_io_to_pes_10_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_32_io_to_mem_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_32_io_to_mem_bits; // @[pe.scala 227:13]
  wire  PENetwork_32_io_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_33_clock; // @[pe.scala 227:13]
  wire  PENetwork_33_io_to_pes_0_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_33_io_to_pes_0_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_33_io_to_pes_0_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_33_io_to_pes_0_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_33_io_to_pes_1_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_33_io_to_pes_1_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_33_io_to_pes_1_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_33_io_to_pes_1_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_33_io_to_pes_1_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_33_io_to_pes_1_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_33_io_to_pes_1_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_33_io_to_pes_2_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_33_io_to_pes_2_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_33_io_to_pes_2_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_33_io_to_pes_2_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_33_io_to_pes_2_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_33_io_to_pes_2_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_33_io_to_pes_2_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_33_io_to_pes_3_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_33_io_to_pes_3_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_33_io_to_pes_3_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_33_io_to_pes_3_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_33_io_to_pes_3_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_33_io_to_pes_3_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_33_io_to_pes_3_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_33_io_to_pes_4_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_33_io_to_pes_4_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_33_io_to_pes_4_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_33_io_to_pes_4_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_33_io_to_pes_4_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_33_io_to_pes_4_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_33_io_to_pes_4_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_33_io_to_pes_5_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_33_io_to_pes_5_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_33_io_to_pes_5_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_33_io_to_pes_5_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_33_io_to_pes_5_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_33_io_to_pes_5_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_33_io_to_pes_5_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_33_io_to_pes_6_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_33_io_to_pes_6_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_33_io_to_pes_6_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_33_io_to_pes_6_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_33_io_to_pes_6_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_33_io_to_pes_6_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_33_io_to_pes_6_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_33_io_to_pes_7_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_33_io_to_pes_7_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_33_io_to_pes_7_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_33_io_to_pes_7_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_33_io_to_pes_7_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_33_io_to_pes_7_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_33_io_to_pes_7_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_33_io_to_pes_8_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_33_io_to_pes_8_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_33_io_to_pes_8_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_33_io_to_pes_8_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_33_io_to_pes_8_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_33_io_to_pes_8_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_33_io_to_pes_8_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_33_io_to_pes_9_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_33_io_to_pes_9_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_33_io_to_pes_9_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_33_io_to_pes_9_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_33_io_to_pes_9_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_33_io_to_pes_9_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_33_io_to_pes_9_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_33_io_to_pes_10_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_33_io_to_pes_10_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_33_io_to_pes_10_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_33_io_to_pes_10_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_33_io_to_pes_10_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_33_io_to_pes_10_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_33_io_to_mem_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_33_io_to_mem_bits; // @[pe.scala 227:13]
  wire  PENetwork_33_io_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_34_clock; // @[pe.scala 227:13]
  wire  PENetwork_34_io_to_pes_0_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_34_io_to_pes_0_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_34_io_to_pes_0_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_34_io_to_pes_0_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_34_io_to_pes_1_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_34_io_to_pes_1_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_34_io_to_pes_1_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_34_io_to_pes_1_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_34_io_to_pes_1_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_34_io_to_pes_1_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_34_io_to_pes_1_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_34_io_to_pes_2_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_34_io_to_pes_2_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_34_io_to_pes_2_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_34_io_to_pes_2_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_34_io_to_pes_2_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_34_io_to_pes_2_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_34_io_to_pes_2_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_34_io_to_pes_3_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_34_io_to_pes_3_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_34_io_to_pes_3_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_34_io_to_pes_3_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_34_io_to_pes_3_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_34_io_to_pes_3_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_34_io_to_pes_3_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_34_io_to_pes_4_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_34_io_to_pes_4_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_34_io_to_pes_4_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_34_io_to_pes_4_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_34_io_to_pes_4_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_34_io_to_pes_4_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_34_io_to_pes_4_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_34_io_to_pes_5_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_34_io_to_pes_5_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_34_io_to_pes_5_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_34_io_to_pes_5_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_34_io_to_pes_5_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_34_io_to_pes_5_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_34_io_to_pes_5_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_34_io_to_pes_6_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_34_io_to_pes_6_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_34_io_to_pes_6_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_34_io_to_pes_6_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_34_io_to_pes_6_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_34_io_to_pes_6_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_34_io_to_pes_6_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_34_io_to_pes_7_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_34_io_to_pes_7_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_34_io_to_pes_7_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_34_io_to_pes_7_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_34_io_to_pes_7_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_34_io_to_pes_7_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_34_io_to_pes_7_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_34_io_to_pes_8_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_34_io_to_pes_8_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_34_io_to_pes_8_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_34_io_to_pes_8_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_34_io_to_pes_8_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_34_io_to_pes_8_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_34_io_to_pes_8_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_34_io_to_pes_9_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_34_io_to_pes_9_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_34_io_to_pes_9_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_34_io_to_pes_9_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_34_io_to_pes_9_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_34_io_to_pes_9_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_34_io_to_pes_9_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_34_io_to_pes_10_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_34_io_to_pes_10_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_34_io_to_pes_10_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_34_io_to_pes_10_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_34_io_to_pes_10_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_34_io_to_pes_10_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_34_io_to_mem_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_34_io_to_mem_bits; // @[pe.scala 227:13]
  wire  PENetwork_34_io_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_35_clock; // @[pe.scala 227:13]
  wire  PENetwork_35_io_to_pes_0_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_35_io_to_pes_0_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_35_io_to_pes_0_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_35_io_to_pes_0_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_35_io_to_pes_1_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_35_io_to_pes_1_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_35_io_to_pes_1_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_35_io_to_pes_1_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_35_io_to_pes_1_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_35_io_to_pes_1_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_35_io_to_pes_1_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_35_io_to_pes_2_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_35_io_to_pes_2_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_35_io_to_pes_2_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_35_io_to_pes_2_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_35_io_to_pes_2_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_35_io_to_pes_2_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_35_io_to_pes_2_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_35_io_to_pes_3_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_35_io_to_pes_3_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_35_io_to_pes_3_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_35_io_to_pes_3_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_35_io_to_pes_3_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_35_io_to_pes_3_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_35_io_to_pes_3_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_35_io_to_pes_4_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_35_io_to_pes_4_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_35_io_to_pes_4_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_35_io_to_pes_4_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_35_io_to_pes_4_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_35_io_to_pes_4_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_35_io_to_pes_4_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_35_io_to_pes_5_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_35_io_to_pes_5_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_35_io_to_pes_5_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_35_io_to_pes_5_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_35_io_to_pes_5_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_35_io_to_pes_5_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_35_io_to_pes_5_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_35_io_to_pes_6_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_35_io_to_pes_6_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_35_io_to_pes_6_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_35_io_to_pes_6_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_35_io_to_pes_6_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_35_io_to_pes_6_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_35_io_to_pes_6_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_35_io_to_pes_7_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_35_io_to_pes_7_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_35_io_to_pes_7_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_35_io_to_pes_7_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_35_io_to_pes_7_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_35_io_to_pes_7_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_35_io_to_pes_7_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_35_io_to_pes_8_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_35_io_to_pes_8_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_35_io_to_pes_8_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_35_io_to_pes_8_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_35_io_to_pes_8_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_35_io_to_pes_8_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_35_io_to_pes_8_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_35_io_to_pes_9_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_35_io_to_pes_9_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_35_io_to_pes_9_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_35_io_to_pes_9_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_35_io_to_pes_9_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_35_io_to_pes_9_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_35_io_to_pes_9_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_35_io_to_pes_10_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_35_io_to_pes_10_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_35_io_to_pes_10_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_35_io_to_pes_10_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_35_io_to_pes_10_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_35_io_to_pes_10_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_35_io_to_mem_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_35_io_to_mem_bits; // @[pe.scala 227:13]
  wire  PENetwork_35_io_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_36_clock; // @[pe.scala 227:13]
  wire  PENetwork_36_io_to_pes_0_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_36_io_to_pes_0_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_36_io_to_pes_0_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_36_io_to_pes_0_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_36_io_to_pes_1_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_36_io_to_pes_1_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_36_io_to_pes_1_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_36_io_to_pes_1_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_36_io_to_pes_1_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_36_io_to_pes_1_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_36_io_to_pes_1_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_36_io_to_pes_2_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_36_io_to_pes_2_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_36_io_to_pes_2_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_36_io_to_pes_2_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_36_io_to_pes_2_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_36_io_to_pes_2_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_36_io_to_pes_2_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_36_io_to_pes_3_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_36_io_to_pes_3_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_36_io_to_pes_3_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_36_io_to_pes_3_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_36_io_to_pes_3_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_36_io_to_pes_3_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_36_io_to_pes_3_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_36_io_to_pes_4_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_36_io_to_pes_4_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_36_io_to_pes_4_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_36_io_to_pes_4_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_36_io_to_pes_4_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_36_io_to_pes_4_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_36_io_to_pes_4_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_36_io_to_pes_5_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_36_io_to_pes_5_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_36_io_to_pes_5_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_36_io_to_pes_5_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_36_io_to_pes_5_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_36_io_to_pes_5_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_36_io_to_pes_5_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_36_io_to_pes_6_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_36_io_to_pes_6_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_36_io_to_pes_6_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_36_io_to_pes_6_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_36_io_to_pes_6_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_36_io_to_pes_6_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_36_io_to_pes_6_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_36_io_to_pes_7_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_36_io_to_pes_7_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_36_io_to_pes_7_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_36_io_to_pes_7_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_36_io_to_pes_7_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_36_io_to_pes_7_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_36_io_to_pes_7_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_36_io_to_pes_8_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_36_io_to_pes_8_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_36_io_to_pes_8_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_36_io_to_pes_8_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_36_io_to_pes_8_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_36_io_to_pes_8_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_36_io_to_pes_8_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_36_io_to_pes_9_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_36_io_to_pes_9_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_36_io_to_pes_9_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_36_io_to_pes_9_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_36_io_to_pes_9_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_36_io_to_pes_9_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_36_io_to_pes_9_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_36_io_to_pes_10_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_36_io_to_pes_10_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_36_io_to_pes_10_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_36_io_to_pes_10_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_36_io_to_pes_10_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_36_io_to_pes_10_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_36_io_to_mem_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_36_io_to_mem_bits; // @[pe.scala 227:13]
  wire  PENetwork_36_io_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_37_clock; // @[pe.scala 227:13]
  wire  PENetwork_37_io_to_pes_0_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_37_io_to_pes_0_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_37_io_to_pes_0_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_37_io_to_pes_0_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_37_io_to_pes_1_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_37_io_to_pes_1_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_37_io_to_pes_1_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_37_io_to_pes_1_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_37_io_to_pes_1_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_37_io_to_pes_1_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_37_io_to_pes_1_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_37_io_to_pes_2_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_37_io_to_pes_2_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_37_io_to_pes_2_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_37_io_to_pes_2_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_37_io_to_pes_2_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_37_io_to_pes_2_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_37_io_to_pes_2_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_37_io_to_pes_3_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_37_io_to_pes_3_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_37_io_to_pes_3_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_37_io_to_pes_3_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_37_io_to_pes_3_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_37_io_to_pes_3_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_37_io_to_pes_3_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_37_io_to_pes_4_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_37_io_to_pes_4_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_37_io_to_pes_4_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_37_io_to_pes_4_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_37_io_to_pes_4_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_37_io_to_pes_4_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_37_io_to_pes_4_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_37_io_to_pes_5_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_37_io_to_pes_5_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_37_io_to_pes_5_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_37_io_to_pes_5_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_37_io_to_pes_5_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_37_io_to_pes_5_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_37_io_to_pes_5_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_37_io_to_pes_6_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_37_io_to_pes_6_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_37_io_to_pes_6_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_37_io_to_pes_6_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_37_io_to_pes_6_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_37_io_to_pes_6_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_37_io_to_pes_6_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_37_io_to_pes_7_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_37_io_to_pes_7_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_37_io_to_pes_7_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_37_io_to_pes_7_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_37_io_to_pes_7_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_37_io_to_pes_7_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_37_io_to_pes_7_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_37_io_to_pes_8_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_37_io_to_pes_8_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_37_io_to_pes_8_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_37_io_to_pes_8_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_37_io_to_pes_8_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_37_io_to_pes_8_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_37_io_to_pes_8_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_37_io_to_pes_9_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_37_io_to_pes_9_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_37_io_to_pes_9_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_37_io_to_pes_9_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_37_io_to_pes_9_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_37_io_to_pes_9_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_37_io_to_pes_9_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_37_io_to_pes_10_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_37_io_to_pes_10_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_37_io_to_pes_10_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_37_io_to_pes_10_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_37_io_to_pes_10_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_37_io_to_pes_10_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_37_io_to_mem_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_37_io_to_mem_bits; // @[pe.scala 227:13]
  wire  PENetwork_37_io_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_38_clock; // @[pe.scala 227:13]
  wire  PENetwork_38_io_to_pes_0_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_38_io_to_pes_0_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_38_io_to_pes_0_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_38_io_to_pes_0_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_38_io_to_pes_1_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_38_io_to_pes_1_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_38_io_to_pes_1_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_38_io_to_pes_1_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_38_io_to_pes_1_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_38_io_to_pes_1_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_38_io_to_pes_1_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_38_io_to_pes_2_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_38_io_to_pes_2_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_38_io_to_pes_2_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_38_io_to_pes_2_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_38_io_to_pes_2_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_38_io_to_pes_2_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_38_io_to_pes_2_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_38_io_to_pes_3_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_38_io_to_pes_3_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_38_io_to_pes_3_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_38_io_to_pes_3_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_38_io_to_pes_3_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_38_io_to_pes_3_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_38_io_to_pes_3_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_38_io_to_pes_4_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_38_io_to_pes_4_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_38_io_to_pes_4_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_38_io_to_pes_4_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_38_io_to_pes_4_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_38_io_to_pes_4_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_38_io_to_pes_4_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_38_io_to_pes_5_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_38_io_to_pes_5_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_38_io_to_pes_5_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_38_io_to_pes_5_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_38_io_to_pes_5_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_38_io_to_pes_5_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_38_io_to_pes_5_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_38_io_to_pes_6_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_38_io_to_pes_6_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_38_io_to_pes_6_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_38_io_to_pes_6_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_38_io_to_pes_6_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_38_io_to_pes_6_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_38_io_to_pes_6_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_38_io_to_pes_7_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_38_io_to_pes_7_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_38_io_to_pes_7_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_38_io_to_pes_7_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_38_io_to_pes_7_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_38_io_to_pes_7_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_38_io_to_pes_7_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_38_io_to_pes_8_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_38_io_to_pes_8_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_38_io_to_pes_8_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_38_io_to_pes_8_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_38_io_to_pes_8_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_38_io_to_pes_8_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_38_io_to_pes_8_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_38_io_to_pes_9_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_38_io_to_pes_9_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_38_io_to_pes_9_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_38_io_to_pes_9_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_38_io_to_pes_9_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_38_io_to_pes_9_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_38_io_to_pes_9_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_38_io_to_pes_10_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_38_io_to_pes_10_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_38_io_to_pes_10_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_38_io_to_pes_10_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_38_io_to_pes_10_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_38_io_to_pes_10_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_38_io_to_mem_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_38_io_to_mem_bits; // @[pe.scala 227:13]
  wire  PENetwork_38_io_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_39_clock; // @[pe.scala 227:13]
  wire  PENetwork_39_io_to_pes_0_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_39_io_to_pes_0_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_39_io_to_pes_0_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_39_io_to_pes_0_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_39_io_to_pes_1_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_39_io_to_pes_1_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_39_io_to_pes_1_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_39_io_to_pes_1_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_39_io_to_pes_1_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_39_io_to_pes_1_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_39_io_to_pes_1_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_39_io_to_pes_2_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_39_io_to_pes_2_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_39_io_to_pes_2_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_39_io_to_pes_2_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_39_io_to_pes_2_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_39_io_to_pes_2_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_39_io_to_pes_2_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_39_io_to_pes_3_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_39_io_to_pes_3_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_39_io_to_pes_3_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_39_io_to_pes_3_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_39_io_to_pes_3_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_39_io_to_pes_3_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_39_io_to_pes_3_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_39_io_to_pes_4_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_39_io_to_pes_4_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_39_io_to_pes_4_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_39_io_to_pes_4_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_39_io_to_pes_4_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_39_io_to_pes_4_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_39_io_to_pes_4_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_39_io_to_pes_5_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_39_io_to_pes_5_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_39_io_to_pes_5_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_39_io_to_pes_5_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_39_io_to_pes_5_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_39_io_to_pes_5_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_39_io_to_pes_5_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_39_io_to_pes_6_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_39_io_to_pes_6_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_39_io_to_pes_6_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_39_io_to_pes_6_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_39_io_to_pes_6_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_39_io_to_pes_6_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_39_io_to_pes_6_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_39_io_to_pes_7_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_39_io_to_pes_7_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_39_io_to_pes_7_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_39_io_to_pes_7_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_39_io_to_pes_7_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_39_io_to_pes_7_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_39_io_to_pes_7_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_39_io_to_pes_8_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_39_io_to_pes_8_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_39_io_to_pes_8_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_39_io_to_pes_8_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_39_io_to_pes_8_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_39_io_to_pes_8_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_39_io_to_pes_8_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_39_io_to_pes_9_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_39_io_to_pes_9_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_39_io_to_pes_9_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_39_io_to_pes_9_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_39_io_to_pes_9_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_39_io_to_pes_9_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_39_io_to_pes_9_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_39_io_to_pes_10_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_39_io_to_pes_10_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_39_io_to_pes_10_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_39_io_to_pes_10_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_39_io_to_pes_10_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_39_io_to_pes_10_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_39_io_to_mem_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_39_io_to_mem_bits; // @[pe.scala 227:13]
  wire  PENetwork_39_io_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_40_clock; // @[pe.scala 227:13]
  wire  PENetwork_40_io_to_pes_0_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_40_io_to_pes_0_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_40_io_to_pes_0_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_40_io_to_pes_0_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_40_io_to_pes_1_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_40_io_to_pes_1_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_40_io_to_pes_1_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_40_io_to_pes_1_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_40_io_to_pes_1_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_40_io_to_pes_1_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_40_io_to_pes_1_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_40_io_to_pes_2_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_40_io_to_pes_2_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_40_io_to_pes_2_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_40_io_to_pes_2_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_40_io_to_pes_2_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_40_io_to_pes_2_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_40_io_to_pes_2_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_40_io_to_pes_3_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_40_io_to_pes_3_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_40_io_to_pes_3_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_40_io_to_pes_3_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_40_io_to_pes_3_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_40_io_to_pes_3_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_40_io_to_pes_3_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_40_io_to_pes_4_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_40_io_to_pes_4_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_40_io_to_pes_4_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_40_io_to_pes_4_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_40_io_to_pes_4_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_40_io_to_pes_4_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_40_io_to_pes_4_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_40_io_to_pes_5_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_40_io_to_pes_5_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_40_io_to_pes_5_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_40_io_to_pes_5_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_40_io_to_pes_5_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_40_io_to_pes_5_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_40_io_to_pes_5_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_40_io_to_pes_6_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_40_io_to_pes_6_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_40_io_to_pes_6_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_40_io_to_pes_6_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_40_io_to_pes_6_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_40_io_to_pes_6_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_40_io_to_pes_6_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_40_io_to_pes_7_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_40_io_to_pes_7_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_40_io_to_pes_7_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_40_io_to_pes_7_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_40_io_to_pes_7_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_40_io_to_pes_7_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_40_io_to_pes_7_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_40_io_to_pes_8_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_40_io_to_pes_8_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_40_io_to_pes_8_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_40_io_to_pes_8_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_40_io_to_pes_8_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_40_io_to_pes_8_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_40_io_to_pes_8_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_40_io_to_pes_9_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_40_io_to_pes_9_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_40_io_to_pes_9_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_40_io_to_pes_9_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_40_io_to_pes_9_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_40_io_to_pes_9_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_40_io_to_pes_9_out_ready; // @[pe.scala 227:13]
  wire  PENetwork_40_io_to_pes_10_in_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_40_io_to_pes_10_in_bits; // @[pe.scala 227:13]
  wire  PENetwork_40_io_to_pes_10_out_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_40_io_to_pes_10_out_bits; // @[pe.scala 227:13]
  wire  PENetwork_40_io_to_pes_10_sig_stat2trans; // @[pe.scala 227:13]
  wire  PENetwork_40_io_to_pes_10_in_ready; // @[pe.scala 227:13]
  wire  PENetwork_40_io_to_mem_valid; // @[pe.scala 227:13]
  wire [255:0] PENetwork_40_io_to_mem_bits; // @[pe.scala 227:13]
  wire  PENetwork_40_io_sig_stat2trans; // @[pe.scala 227:13]
  wire  MemController_clock; // @[pe.scala 306:15]
  wire  MemController_reset; // @[pe.scala 306:15]
  wire  MemController_io_rd_valid; // @[pe.scala 306:15]
  wire  MemController_io_wr_valid; // @[pe.scala 306:15]
  wire  MemController_io_rd_data_valid; // @[pe.scala 306:15]
  wire [31:0] MemController_io_rd_data_bits; // @[pe.scala 306:15]
  wire  MemController_io_wr_data_valid; // @[pe.scala 306:15]
  wire [31:0] MemController_io_wr_data_bits; // @[pe.scala 306:15]
  wire  MemController_1_clock; // @[pe.scala 306:15]
  wire  MemController_1_reset; // @[pe.scala 306:15]
  wire  MemController_1_io_rd_valid; // @[pe.scala 306:15]
  wire  MemController_1_io_wr_valid; // @[pe.scala 306:15]
  wire  MemController_1_io_rd_data_valid; // @[pe.scala 306:15]
  wire [31:0] MemController_1_io_rd_data_bits; // @[pe.scala 306:15]
  wire  MemController_1_io_wr_data_valid; // @[pe.scala 306:15]
  wire [31:0] MemController_1_io_wr_data_bits; // @[pe.scala 306:15]
  wire  MemController_2_clock; // @[pe.scala 306:15]
  wire  MemController_2_reset; // @[pe.scala 306:15]
  wire  MemController_2_io_rd_valid; // @[pe.scala 306:15]
  wire  MemController_2_io_wr_valid; // @[pe.scala 306:15]
  wire  MemController_2_io_rd_data_valid; // @[pe.scala 306:15]
  wire [31:0] MemController_2_io_rd_data_bits; // @[pe.scala 306:15]
  wire  MemController_2_io_wr_data_valid; // @[pe.scala 306:15]
  wire [31:0] MemController_2_io_wr_data_bits; // @[pe.scala 306:15]
  wire  MemController_3_clock; // @[pe.scala 306:15]
  wire  MemController_3_reset; // @[pe.scala 306:15]
  wire  MemController_3_io_rd_valid; // @[pe.scala 306:15]
  wire  MemController_3_io_wr_valid; // @[pe.scala 306:15]
  wire  MemController_3_io_rd_data_valid; // @[pe.scala 306:15]
  wire [31:0] MemController_3_io_rd_data_bits; // @[pe.scala 306:15]
  wire  MemController_3_io_wr_data_valid; // @[pe.scala 306:15]
  wire [31:0] MemController_3_io_wr_data_bits; // @[pe.scala 306:15]
  wire  MemController_4_clock; // @[pe.scala 306:15]
  wire  MemController_4_reset; // @[pe.scala 306:15]
  wire  MemController_4_io_rd_valid; // @[pe.scala 306:15]
  wire  MemController_4_io_wr_valid; // @[pe.scala 306:15]
  wire  MemController_4_io_rd_data_valid; // @[pe.scala 306:15]
  wire [31:0] MemController_4_io_rd_data_bits; // @[pe.scala 306:15]
  wire  MemController_4_io_wr_data_valid; // @[pe.scala 306:15]
  wire [31:0] MemController_4_io_wr_data_bits; // @[pe.scala 306:15]
  wire  MemController_5_clock; // @[pe.scala 306:15]
  wire  MemController_5_reset; // @[pe.scala 306:15]
  wire  MemController_5_io_rd_valid; // @[pe.scala 306:15]
  wire  MemController_5_io_wr_valid; // @[pe.scala 306:15]
  wire  MemController_5_io_rd_data_valid; // @[pe.scala 306:15]
  wire [31:0] MemController_5_io_rd_data_bits; // @[pe.scala 306:15]
  wire  MemController_5_io_wr_data_valid; // @[pe.scala 306:15]
  wire [31:0] MemController_5_io_wr_data_bits; // @[pe.scala 306:15]
  wire  MemController_6_clock; // @[pe.scala 306:15]
  wire  MemController_6_reset; // @[pe.scala 306:15]
  wire  MemController_6_io_rd_valid; // @[pe.scala 306:15]
  wire  MemController_6_io_wr_valid; // @[pe.scala 306:15]
  wire  MemController_6_io_rd_data_valid; // @[pe.scala 306:15]
  wire [31:0] MemController_6_io_rd_data_bits; // @[pe.scala 306:15]
  wire  MemController_6_io_wr_data_valid; // @[pe.scala 306:15]
  wire [31:0] MemController_6_io_wr_data_bits; // @[pe.scala 306:15]
  wire  MemController_7_clock; // @[pe.scala 306:15]
  wire  MemController_7_reset; // @[pe.scala 306:15]
  wire  MemController_7_io_rd_valid; // @[pe.scala 306:15]
  wire  MemController_7_io_wr_valid; // @[pe.scala 306:15]
  wire  MemController_7_io_rd_data_valid; // @[pe.scala 306:15]
  wire [31:0] MemController_7_io_rd_data_bits; // @[pe.scala 306:15]
  wire  MemController_7_io_wr_data_valid; // @[pe.scala 306:15]
  wire [31:0] MemController_7_io_wr_data_bits; // @[pe.scala 306:15]
  wire  MemController_8_clock; // @[pe.scala 306:15]
  wire  MemController_8_reset; // @[pe.scala 306:15]
  wire  MemController_8_io_rd_valid; // @[pe.scala 306:15]
  wire  MemController_8_io_wr_valid; // @[pe.scala 306:15]
  wire  MemController_8_io_rd_data_valid; // @[pe.scala 306:15]
  wire [31:0] MemController_8_io_rd_data_bits; // @[pe.scala 306:15]
  wire  MemController_8_io_wr_data_valid; // @[pe.scala 306:15]
  wire [31:0] MemController_8_io_wr_data_bits; // @[pe.scala 306:15]
  wire  MemController_9_clock; // @[pe.scala 306:15]
  wire  MemController_9_reset; // @[pe.scala 306:15]
  wire  MemController_9_io_rd_valid; // @[pe.scala 306:15]
  wire  MemController_9_io_wr_valid; // @[pe.scala 306:15]
  wire  MemController_9_io_rd_data_valid; // @[pe.scala 306:15]
  wire [31:0] MemController_9_io_rd_data_bits; // @[pe.scala 306:15]
  wire  MemController_9_io_wr_data_valid; // @[pe.scala 306:15]
  wire [31:0] MemController_9_io_wr_data_bits; // @[pe.scala 306:15]
  wire  MemController_10_clock; // @[pe.scala 306:15]
  wire  MemController_10_reset; // @[pe.scala 306:15]
  wire  MemController_10_io_rd_valid; // @[pe.scala 306:15]
  wire  MemController_10_io_wr_valid; // @[pe.scala 306:15]
  wire  MemController_10_io_rd_data_valid; // @[pe.scala 306:15]
  wire [31:0] MemController_10_io_rd_data_bits; // @[pe.scala 306:15]
  wire  MemController_10_io_wr_data_valid; // @[pe.scala 306:15]
  wire [31:0] MemController_10_io_wr_data_bits; // @[pe.scala 306:15]
  wire  MemController_11_clock; // @[pe.scala 306:15]
  wire  MemController_11_reset; // @[pe.scala 306:15]
  wire  MemController_11_io_rd_valid; // @[pe.scala 306:15]
  wire  MemController_11_io_wr_valid; // @[pe.scala 306:15]
  wire  MemController_11_io_rd_data_valid; // @[pe.scala 306:15]
  wire [255:0] MemController_11_io_rd_data_bits; // @[pe.scala 306:15]
  wire  MemController_11_io_wr_data_valid; // @[pe.scala 306:15]
  wire [255:0] MemController_11_io_wr_data_bits; // @[pe.scala 306:15]
  wire  MemController_12_clock; // @[pe.scala 306:15]
  wire  MemController_12_reset; // @[pe.scala 306:15]
  wire  MemController_12_io_rd_valid; // @[pe.scala 306:15]
  wire  MemController_12_io_wr_valid; // @[pe.scala 306:15]
  wire  MemController_12_io_rd_data_valid; // @[pe.scala 306:15]
  wire [255:0] MemController_12_io_rd_data_bits; // @[pe.scala 306:15]
  wire  MemController_12_io_wr_data_valid; // @[pe.scala 306:15]
  wire [255:0] MemController_12_io_wr_data_bits; // @[pe.scala 306:15]
  wire  MemController_13_clock; // @[pe.scala 306:15]
  wire  MemController_13_reset; // @[pe.scala 306:15]
  wire  MemController_13_io_rd_valid; // @[pe.scala 306:15]
  wire  MemController_13_io_wr_valid; // @[pe.scala 306:15]
  wire  MemController_13_io_rd_data_valid; // @[pe.scala 306:15]
  wire [255:0] MemController_13_io_rd_data_bits; // @[pe.scala 306:15]
  wire  MemController_13_io_wr_data_valid; // @[pe.scala 306:15]
  wire [255:0] MemController_13_io_wr_data_bits; // @[pe.scala 306:15]
  wire  MemController_14_clock; // @[pe.scala 306:15]
  wire  MemController_14_reset; // @[pe.scala 306:15]
  wire  MemController_14_io_rd_valid; // @[pe.scala 306:15]
  wire  MemController_14_io_wr_valid; // @[pe.scala 306:15]
  wire  MemController_14_io_rd_data_valid; // @[pe.scala 306:15]
  wire [255:0] MemController_14_io_rd_data_bits; // @[pe.scala 306:15]
  wire  MemController_14_io_wr_data_valid; // @[pe.scala 306:15]
  wire [255:0] MemController_14_io_wr_data_bits; // @[pe.scala 306:15]
  wire  MemController_15_clock; // @[pe.scala 306:15]
  wire  MemController_15_reset; // @[pe.scala 306:15]
  wire  MemController_15_io_rd_valid; // @[pe.scala 306:15]
  wire  MemController_15_io_wr_valid; // @[pe.scala 306:15]
  wire  MemController_15_io_rd_data_valid; // @[pe.scala 306:15]
  wire [255:0] MemController_15_io_rd_data_bits; // @[pe.scala 306:15]
  wire  MemController_15_io_wr_data_valid; // @[pe.scala 306:15]
  wire [255:0] MemController_15_io_wr_data_bits; // @[pe.scala 306:15]
  wire  MemController_16_clock; // @[pe.scala 306:15]
  wire  MemController_16_reset; // @[pe.scala 306:15]
  wire  MemController_16_io_rd_valid; // @[pe.scala 306:15]
  wire  MemController_16_io_wr_valid; // @[pe.scala 306:15]
  wire  MemController_16_io_rd_data_valid; // @[pe.scala 306:15]
  wire [255:0] MemController_16_io_rd_data_bits; // @[pe.scala 306:15]
  wire  MemController_16_io_wr_data_valid; // @[pe.scala 306:15]
  wire [255:0] MemController_16_io_wr_data_bits; // @[pe.scala 306:15]
  wire  MemController_17_clock; // @[pe.scala 306:15]
  wire  MemController_17_reset; // @[pe.scala 306:15]
  wire  MemController_17_io_rd_valid; // @[pe.scala 306:15]
  wire  MemController_17_io_wr_valid; // @[pe.scala 306:15]
  wire  MemController_17_io_rd_data_valid; // @[pe.scala 306:15]
  wire [255:0] MemController_17_io_rd_data_bits; // @[pe.scala 306:15]
  wire  MemController_17_io_wr_data_valid; // @[pe.scala 306:15]
  wire [255:0] MemController_17_io_wr_data_bits; // @[pe.scala 306:15]
  wire  MemController_18_clock; // @[pe.scala 306:15]
  wire  MemController_18_reset; // @[pe.scala 306:15]
  wire  MemController_18_io_rd_valid; // @[pe.scala 306:15]
  wire  MemController_18_io_wr_valid; // @[pe.scala 306:15]
  wire  MemController_18_io_rd_data_valid; // @[pe.scala 306:15]
  wire [255:0] MemController_18_io_rd_data_bits; // @[pe.scala 306:15]
  wire  MemController_18_io_wr_data_valid; // @[pe.scala 306:15]
  wire [255:0] MemController_18_io_wr_data_bits; // @[pe.scala 306:15]
  wire  MemController_19_clock; // @[pe.scala 306:15]
  wire  MemController_19_reset; // @[pe.scala 306:15]
  wire  MemController_19_io_rd_valid; // @[pe.scala 306:15]
  wire  MemController_19_io_wr_valid; // @[pe.scala 306:15]
  wire  MemController_19_io_rd_data_valid; // @[pe.scala 306:15]
  wire [255:0] MemController_19_io_rd_data_bits; // @[pe.scala 306:15]
  wire  MemController_19_io_wr_data_valid; // @[pe.scala 306:15]
  wire [255:0] MemController_19_io_wr_data_bits; // @[pe.scala 306:15]
  wire  MemController_20_clock; // @[pe.scala 306:15]
  wire  MemController_20_reset; // @[pe.scala 306:15]
  wire  MemController_20_io_rd_valid; // @[pe.scala 306:15]
  wire  MemController_20_io_wr_valid; // @[pe.scala 306:15]
  wire  MemController_20_io_rd_data_valid; // @[pe.scala 306:15]
  wire [255:0] MemController_20_io_rd_data_bits; // @[pe.scala 306:15]
  wire  MemController_20_io_wr_data_valid; // @[pe.scala 306:15]
  wire [255:0] MemController_20_io_wr_data_bits; // @[pe.scala 306:15]
  wire  MemController_21_clock; // @[pe.scala 306:15]
  wire  MemController_21_reset; // @[pe.scala 306:15]
  wire  MemController_21_io_rd_valid; // @[pe.scala 306:15]
  wire  MemController_21_io_wr_valid; // @[pe.scala 306:15]
  wire  MemController_21_io_rd_data_valid; // @[pe.scala 306:15]
  wire [255:0] MemController_21_io_rd_data_bits; // @[pe.scala 306:15]
  wire  MemController_21_io_wr_data_valid; // @[pe.scala 306:15]
  wire [255:0] MemController_21_io_wr_data_bits; // @[pe.scala 306:15]
  wire  MemController_22_clock; // @[pe.scala 306:15]
  wire  MemController_22_reset; // @[pe.scala 306:15]
  wire  MemController_22_io_rd_valid; // @[pe.scala 306:15]
  wire  MemController_22_io_wr_valid; // @[pe.scala 306:15]
  wire  MemController_22_io_rd_data_valid; // @[pe.scala 306:15]
  wire [255:0] MemController_22_io_rd_data_bits; // @[pe.scala 306:15]
  wire  MemController_22_io_wr_data_valid; // @[pe.scala 306:15]
  wire [255:0] MemController_22_io_wr_data_bits; // @[pe.scala 306:15]
  wire  MemController_23_clock; // @[pe.scala 306:15]
  wire  MemController_23_reset; // @[pe.scala 306:15]
  wire  MemController_23_io_rd_valid; // @[pe.scala 306:15]
  wire  MemController_23_io_wr_valid; // @[pe.scala 306:15]
  wire  MemController_23_io_rd_data_valid; // @[pe.scala 306:15]
  wire [255:0] MemController_23_io_rd_data_bits; // @[pe.scala 306:15]
  wire  MemController_23_io_wr_data_valid; // @[pe.scala 306:15]
  wire [255:0] MemController_23_io_wr_data_bits; // @[pe.scala 306:15]
  wire  MemController_24_clock; // @[pe.scala 306:15]
  wire  MemController_24_reset; // @[pe.scala 306:15]
  wire  MemController_24_io_rd_valid; // @[pe.scala 306:15]
  wire  MemController_24_io_wr_valid; // @[pe.scala 306:15]
  wire  MemController_24_io_rd_data_valid; // @[pe.scala 306:15]
  wire [255:0] MemController_24_io_rd_data_bits; // @[pe.scala 306:15]
  wire  MemController_24_io_wr_data_valid; // @[pe.scala 306:15]
  wire [255:0] MemController_24_io_wr_data_bits; // @[pe.scala 306:15]
  wire  MemController_25_clock; // @[pe.scala 306:15]
  wire  MemController_25_reset; // @[pe.scala 306:15]
  wire  MemController_25_io_rd_valid; // @[pe.scala 306:15]
  wire  MemController_25_io_wr_valid; // @[pe.scala 306:15]
  wire  MemController_25_io_rd_data_valid; // @[pe.scala 306:15]
  wire [255:0] MemController_25_io_rd_data_bits; // @[pe.scala 306:15]
  wire  MemController_25_io_wr_data_valid; // @[pe.scala 306:15]
  wire [255:0] MemController_25_io_wr_data_bits; // @[pe.scala 306:15]
  wire  MemController_26_clock; // @[pe.scala 304:15]
  wire  MemController_26_reset; // @[pe.scala 304:15]
  wire  MemController_26_io_rd_valid; // @[pe.scala 304:15]
  wire  MemController_26_io_wr_valid; // @[pe.scala 304:15]
  wire  MemController_26_io_rd_data_valid; // @[pe.scala 304:15]
  wire [255:0] MemController_26_io_rd_data_bits; // @[pe.scala 304:15]
  wire  MemController_26_io_wr_data_valid; // @[pe.scala 304:15]
  wire [255:0] MemController_26_io_wr_data_bits; // @[pe.scala 304:15]
  wire  MemController_27_clock; // @[pe.scala 304:15]
  wire  MemController_27_reset; // @[pe.scala 304:15]
  wire  MemController_27_io_rd_valid; // @[pe.scala 304:15]
  wire  MemController_27_io_wr_valid; // @[pe.scala 304:15]
  wire  MemController_27_io_rd_data_valid; // @[pe.scala 304:15]
  wire [255:0] MemController_27_io_rd_data_bits; // @[pe.scala 304:15]
  wire  MemController_27_io_wr_data_valid; // @[pe.scala 304:15]
  wire [255:0] MemController_27_io_wr_data_bits; // @[pe.scala 304:15]
  wire  MemController_28_clock; // @[pe.scala 304:15]
  wire  MemController_28_reset; // @[pe.scala 304:15]
  wire  MemController_28_io_rd_valid; // @[pe.scala 304:15]
  wire  MemController_28_io_wr_valid; // @[pe.scala 304:15]
  wire  MemController_28_io_rd_data_valid; // @[pe.scala 304:15]
  wire [255:0] MemController_28_io_rd_data_bits; // @[pe.scala 304:15]
  wire  MemController_28_io_wr_data_valid; // @[pe.scala 304:15]
  wire [255:0] MemController_28_io_wr_data_bits; // @[pe.scala 304:15]
  wire  MemController_29_clock; // @[pe.scala 304:15]
  wire  MemController_29_reset; // @[pe.scala 304:15]
  wire  MemController_29_io_rd_valid; // @[pe.scala 304:15]
  wire  MemController_29_io_wr_valid; // @[pe.scala 304:15]
  wire  MemController_29_io_rd_data_valid; // @[pe.scala 304:15]
  wire [255:0] MemController_29_io_rd_data_bits; // @[pe.scala 304:15]
  wire  MemController_29_io_wr_data_valid; // @[pe.scala 304:15]
  wire [255:0] MemController_29_io_wr_data_bits; // @[pe.scala 304:15]
  wire  MemController_30_clock; // @[pe.scala 304:15]
  wire  MemController_30_reset; // @[pe.scala 304:15]
  wire  MemController_30_io_rd_valid; // @[pe.scala 304:15]
  wire  MemController_30_io_wr_valid; // @[pe.scala 304:15]
  wire  MemController_30_io_rd_data_valid; // @[pe.scala 304:15]
  wire [255:0] MemController_30_io_rd_data_bits; // @[pe.scala 304:15]
  wire  MemController_30_io_wr_data_valid; // @[pe.scala 304:15]
  wire [255:0] MemController_30_io_wr_data_bits; // @[pe.scala 304:15]
  wire  MemController_31_clock; // @[pe.scala 304:15]
  wire  MemController_31_reset; // @[pe.scala 304:15]
  wire  MemController_31_io_rd_valid; // @[pe.scala 304:15]
  wire  MemController_31_io_wr_valid; // @[pe.scala 304:15]
  wire  MemController_31_io_rd_data_valid; // @[pe.scala 304:15]
  wire [255:0] MemController_31_io_rd_data_bits; // @[pe.scala 304:15]
  wire  MemController_31_io_wr_data_valid; // @[pe.scala 304:15]
  wire [255:0] MemController_31_io_wr_data_bits; // @[pe.scala 304:15]
  wire  MemController_32_clock; // @[pe.scala 304:15]
  wire  MemController_32_reset; // @[pe.scala 304:15]
  wire  MemController_32_io_rd_valid; // @[pe.scala 304:15]
  wire  MemController_32_io_wr_valid; // @[pe.scala 304:15]
  wire  MemController_32_io_rd_data_valid; // @[pe.scala 304:15]
  wire [255:0] MemController_32_io_rd_data_bits; // @[pe.scala 304:15]
  wire  MemController_32_io_wr_data_valid; // @[pe.scala 304:15]
  wire [255:0] MemController_32_io_wr_data_bits; // @[pe.scala 304:15]
  wire  MemController_33_clock; // @[pe.scala 304:15]
  wire  MemController_33_reset; // @[pe.scala 304:15]
  wire  MemController_33_io_rd_valid; // @[pe.scala 304:15]
  wire  MemController_33_io_wr_valid; // @[pe.scala 304:15]
  wire  MemController_33_io_rd_data_valid; // @[pe.scala 304:15]
  wire [255:0] MemController_33_io_rd_data_bits; // @[pe.scala 304:15]
  wire  MemController_33_io_wr_data_valid; // @[pe.scala 304:15]
  wire [255:0] MemController_33_io_wr_data_bits; // @[pe.scala 304:15]
  wire  MemController_34_clock; // @[pe.scala 304:15]
  wire  MemController_34_reset; // @[pe.scala 304:15]
  wire  MemController_34_io_rd_valid; // @[pe.scala 304:15]
  wire  MemController_34_io_wr_valid; // @[pe.scala 304:15]
  wire  MemController_34_io_rd_data_valid; // @[pe.scala 304:15]
  wire [255:0] MemController_34_io_rd_data_bits; // @[pe.scala 304:15]
  wire  MemController_34_io_wr_data_valid; // @[pe.scala 304:15]
  wire [255:0] MemController_34_io_wr_data_bits; // @[pe.scala 304:15]
  wire  MemController_35_clock; // @[pe.scala 304:15]
  wire  MemController_35_reset; // @[pe.scala 304:15]
  wire  MemController_35_io_rd_valid; // @[pe.scala 304:15]
  wire  MemController_35_io_wr_valid; // @[pe.scala 304:15]
  wire  MemController_35_io_rd_data_valid; // @[pe.scala 304:15]
  wire [255:0] MemController_35_io_rd_data_bits; // @[pe.scala 304:15]
  wire  MemController_35_io_wr_data_valid; // @[pe.scala 304:15]
  wire [255:0] MemController_35_io_wr_data_bits; // @[pe.scala 304:15]
  wire  MemController_36_clock; // @[pe.scala 304:15]
  wire  MemController_36_reset; // @[pe.scala 304:15]
  wire  MemController_36_io_rd_valid; // @[pe.scala 304:15]
  wire  MemController_36_io_wr_valid; // @[pe.scala 304:15]
  wire  MemController_36_io_rd_data_valid; // @[pe.scala 304:15]
  wire [255:0] MemController_36_io_rd_data_bits; // @[pe.scala 304:15]
  wire  MemController_36_io_wr_data_valid; // @[pe.scala 304:15]
  wire [255:0] MemController_36_io_wr_data_bits; // @[pe.scala 304:15]
  wire  MemController_37_clock; // @[pe.scala 304:15]
  wire  MemController_37_reset; // @[pe.scala 304:15]
  wire  MemController_37_io_rd_valid; // @[pe.scala 304:15]
  wire  MemController_37_io_wr_valid; // @[pe.scala 304:15]
  wire  MemController_37_io_rd_data_valid; // @[pe.scala 304:15]
  wire [255:0] MemController_37_io_rd_data_bits; // @[pe.scala 304:15]
  wire  MemController_37_io_wr_data_valid; // @[pe.scala 304:15]
  wire [255:0] MemController_37_io_wr_data_bits; // @[pe.scala 304:15]
  wire  MemController_38_clock; // @[pe.scala 304:15]
  wire  MemController_38_reset; // @[pe.scala 304:15]
  wire  MemController_38_io_rd_valid; // @[pe.scala 304:15]
  wire  MemController_38_io_wr_valid; // @[pe.scala 304:15]
  wire  MemController_38_io_rd_data_valid; // @[pe.scala 304:15]
  wire [255:0] MemController_38_io_rd_data_bits; // @[pe.scala 304:15]
  wire  MemController_38_io_wr_data_valid; // @[pe.scala 304:15]
  wire [255:0] MemController_38_io_wr_data_bits; // @[pe.scala 304:15]
  wire  MemController_39_clock; // @[pe.scala 304:15]
  wire  MemController_39_reset; // @[pe.scala 304:15]
  wire  MemController_39_io_rd_valid; // @[pe.scala 304:15]
  wire  MemController_39_io_wr_valid; // @[pe.scala 304:15]
  wire  MemController_39_io_rd_data_valid; // @[pe.scala 304:15]
  wire [255:0] MemController_39_io_rd_data_bits; // @[pe.scala 304:15]
  wire  MemController_39_io_wr_data_valid; // @[pe.scala 304:15]
  wire [255:0] MemController_39_io_wr_data_bits; // @[pe.scala 304:15]
  wire  MemController_40_clock; // @[pe.scala 304:15]
  wire  MemController_40_reset; // @[pe.scala 304:15]
  wire  MemController_40_io_rd_valid; // @[pe.scala 304:15]
  wire  MemController_40_io_wr_valid; // @[pe.scala 304:15]
  wire  MemController_40_io_rd_data_valid; // @[pe.scala 304:15]
  wire [255:0] MemController_40_io_rd_data_bits; // @[pe.scala 304:15]
  wire  MemController_40_io_wr_data_valid; // @[pe.scala 304:15]
  wire [255:0] MemController_40_io_wr_data_bits; // @[pe.scala 304:15]
  wire  _T_1 = ~reset; // @[pe.scala 163:9]
  MultiDimTime MultiDimTime ( // @[pe.scala 162:25]
    .clock(MultiDimTime_clock),
    .reset(MultiDimTime_reset),
    .io_in(MultiDimTime_io_in),
    .io_out_0(MultiDimTime_io_out_0),
    .io_out_1(MultiDimTime_io_out_1),
    .io_out_2(MultiDimTime_io_out_2),
    .io_index_0(MultiDimTime_io_index_0),
    .io_index_1(MultiDimTime_io_index_1),
    .io_index_2(MultiDimTime_io_index_2)
  );
  PE PE ( // @[pe.scala 184:13]
    .clock(PE_clock),
    .reset(PE_reset),
    .io_data_2_in_valid(PE_io_data_2_in_valid),
    .io_data_2_in_bits(PE_io_data_2_in_bits),
    .io_data_2_out_valid(PE_io_data_2_out_valid),
    .io_data_2_out_bits(PE_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_io_data_2_in_ready),
    .io_data_2_out_ready(PE_io_data_2_out_ready),
    .io_data_1_in_valid(PE_io_data_1_in_valid),
    .io_data_1_in_bits(PE_io_data_1_in_bits),
    .io_data_1_out_valid(PE_io_data_1_out_valid),
    .io_data_1_out_bits(PE_io_data_1_out_bits),
    .io_data_0_in_valid(PE_io_data_0_in_valid),
    .io_data_0_in_bits(PE_io_data_0_in_bits),
    .io_data_0_out_valid(PE_io_data_0_out_valid),
    .io_data_0_out_bits(PE_io_data_0_out_bits)
  );
  PE PE_1 ( // @[pe.scala 184:13]
    .clock(PE_1_clock),
    .reset(PE_1_reset),
    .io_data_2_in_valid(PE_1_io_data_2_in_valid),
    .io_data_2_in_bits(PE_1_io_data_2_in_bits),
    .io_data_2_out_valid(PE_1_io_data_2_out_valid),
    .io_data_2_out_bits(PE_1_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_1_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_1_io_data_2_in_ready),
    .io_data_2_out_ready(PE_1_io_data_2_out_ready),
    .io_data_1_in_valid(PE_1_io_data_1_in_valid),
    .io_data_1_in_bits(PE_1_io_data_1_in_bits),
    .io_data_1_out_valid(PE_1_io_data_1_out_valid),
    .io_data_1_out_bits(PE_1_io_data_1_out_bits),
    .io_data_0_in_valid(PE_1_io_data_0_in_valid),
    .io_data_0_in_bits(PE_1_io_data_0_in_bits),
    .io_data_0_out_valid(PE_1_io_data_0_out_valid),
    .io_data_0_out_bits(PE_1_io_data_0_out_bits)
  );
  PE PE_2 ( // @[pe.scala 184:13]
    .clock(PE_2_clock),
    .reset(PE_2_reset),
    .io_data_2_in_valid(PE_2_io_data_2_in_valid),
    .io_data_2_in_bits(PE_2_io_data_2_in_bits),
    .io_data_2_out_valid(PE_2_io_data_2_out_valid),
    .io_data_2_out_bits(PE_2_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_2_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_2_io_data_2_in_ready),
    .io_data_2_out_ready(PE_2_io_data_2_out_ready),
    .io_data_1_in_valid(PE_2_io_data_1_in_valid),
    .io_data_1_in_bits(PE_2_io_data_1_in_bits),
    .io_data_1_out_valid(PE_2_io_data_1_out_valid),
    .io_data_1_out_bits(PE_2_io_data_1_out_bits),
    .io_data_0_in_valid(PE_2_io_data_0_in_valid),
    .io_data_0_in_bits(PE_2_io_data_0_in_bits),
    .io_data_0_out_valid(PE_2_io_data_0_out_valid),
    .io_data_0_out_bits(PE_2_io_data_0_out_bits)
  );
  PE PE_3 ( // @[pe.scala 184:13]
    .clock(PE_3_clock),
    .reset(PE_3_reset),
    .io_data_2_in_valid(PE_3_io_data_2_in_valid),
    .io_data_2_in_bits(PE_3_io_data_2_in_bits),
    .io_data_2_out_valid(PE_3_io_data_2_out_valid),
    .io_data_2_out_bits(PE_3_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_3_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_3_io_data_2_in_ready),
    .io_data_2_out_ready(PE_3_io_data_2_out_ready),
    .io_data_1_in_valid(PE_3_io_data_1_in_valid),
    .io_data_1_in_bits(PE_3_io_data_1_in_bits),
    .io_data_1_out_valid(PE_3_io_data_1_out_valid),
    .io_data_1_out_bits(PE_3_io_data_1_out_bits),
    .io_data_0_in_valid(PE_3_io_data_0_in_valid),
    .io_data_0_in_bits(PE_3_io_data_0_in_bits),
    .io_data_0_out_valid(PE_3_io_data_0_out_valid),
    .io_data_0_out_bits(PE_3_io_data_0_out_bits)
  );
  PE PE_4 ( // @[pe.scala 184:13]
    .clock(PE_4_clock),
    .reset(PE_4_reset),
    .io_data_2_in_valid(PE_4_io_data_2_in_valid),
    .io_data_2_in_bits(PE_4_io_data_2_in_bits),
    .io_data_2_out_valid(PE_4_io_data_2_out_valid),
    .io_data_2_out_bits(PE_4_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_4_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_4_io_data_2_in_ready),
    .io_data_2_out_ready(PE_4_io_data_2_out_ready),
    .io_data_1_in_valid(PE_4_io_data_1_in_valid),
    .io_data_1_in_bits(PE_4_io_data_1_in_bits),
    .io_data_1_out_valid(PE_4_io_data_1_out_valid),
    .io_data_1_out_bits(PE_4_io_data_1_out_bits),
    .io_data_0_in_valid(PE_4_io_data_0_in_valid),
    .io_data_0_in_bits(PE_4_io_data_0_in_bits),
    .io_data_0_out_valid(PE_4_io_data_0_out_valid),
    .io_data_0_out_bits(PE_4_io_data_0_out_bits)
  );
  PE PE_5 ( // @[pe.scala 184:13]
    .clock(PE_5_clock),
    .reset(PE_5_reset),
    .io_data_2_in_valid(PE_5_io_data_2_in_valid),
    .io_data_2_in_bits(PE_5_io_data_2_in_bits),
    .io_data_2_out_valid(PE_5_io_data_2_out_valid),
    .io_data_2_out_bits(PE_5_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_5_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_5_io_data_2_in_ready),
    .io_data_2_out_ready(PE_5_io_data_2_out_ready),
    .io_data_1_in_valid(PE_5_io_data_1_in_valid),
    .io_data_1_in_bits(PE_5_io_data_1_in_bits),
    .io_data_1_out_valid(PE_5_io_data_1_out_valid),
    .io_data_1_out_bits(PE_5_io_data_1_out_bits),
    .io_data_0_in_valid(PE_5_io_data_0_in_valid),
    .io_data_0_in_bits(PE_5_io_data_0_in_bits),
    .io_data_0_out_valid(PE_5_io_data_0_out_valid),
    .io_data_0_out_bits(PE_5_io_data_0_out_bits)
  );
  PE PE_6 ( // @[pe.scala 184:13]
    .clock(PE_6_clock),
    .reset(PE_6_reset),
    .io_data_2_in_valid(PE_6_io_data_2_in_valid),
    .io_data_2_in_bits(PE_6_io_data_2_in_bits),
    .io_data_2_out_valid(PE_6_io_data_2_out_valid),
    .io_data_2_out_bits(PE_6_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_6_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_6_io_data_2_in_ready),
    .io_data_2_out_ready(PE_6_io_data_2_out_ready),
    .io_data_1_in_valid(PE_6_io_data_1_in_valid),
    .io_data_1_in_bits(PE_6_io_data_1_in_bits),
    .io_data_1_out_valid(PE_6_io_data_1_out_valid),
    .io_data_1_out_bits(PE_6_io_data_1_out_bits),
    .io_data_0_in_valid(PE_6_io_data_0_in_valid),
    .io_data_0_in_bits(PE_6_io_data_0_in_bits),
    .io_data_0_out_valid(PE_6_io_data_0_out_valid),
    .io_data_0_out_bits(PE_6_io_data_0_out_bits)
  );
  PE PE_7 ( // @[pe.scala 184:13]
    .clock(PE_7_clock),
    .reset(PE_7_reset),
    .io_data_2_in_valid(PE_7_io_data_2_in_valid),
    .io_data_2_in_bits(PE_7_io_data_2_in_bits),
    .io_data_2_out_valid(PE_7_io_data_2_out_valid),
    .io_data_2_out_bits(PE_7_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_7_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_7_io_data_2_in_ready),
    .io_data_2_out_ready(PE_7_io_data_2_out_ready),
    .io_data_1_in_valid(PE_7_io_data_1_in_valid),
    .io_data_1_in_bits(PE_7_io_data_1_in_bits),
    .io_data_1_out_valid(PE_7_io_data_1_out_valid),
    .io_data_1_out_bits(PE_7_io_data_1_out_bits),
    .io_data_0_in_valid(PE_7_io_data_0_in_valid),
    .io_data_0_in_bits(PE_7_io_data_0_in_bits),
    .io_data_0_out_valid(PE_7_io_data_0_out_valid),
    .io_data_0_out_bits(PE_7_io_data_0_out_bits)
  );
  PE PE_8 ( // @[pe.scala 184:13]
    .clock(PE_8_clock),
    .reset(PE_8_reset),
    .io_data_2_in_valid(PE_8_io_data_2_in_valid),
    .io_data_2_in_bits(PE_8_io_data_2_in_bits),
    .io_data_2_out_valid(PE_8_io_data_2_out_valid),
    .io_data_2_out_bits(PE_8_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_8_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_8_io_data_2_in_ready),
    .io_data_2_out_ready(PE_8_io_data_2_out_ready),
    .io_data_1_in_valid(PE_8_io_data_1_in_valid),
    .io_data_1_in_bits(PE_8_io_data_1_in_bits),
    .io_data_1_out_valid(PE_8_io_data_1_out_valid),
    .io_data_1_out_bits(PE_8_io_data_1_out_bits),
    .io_data_0_in_valid(PE_8_io_data_0_in_valid),
    .io_data_0_in_bits(PE_8_io_data_0_in_bits),
    .io_data_0_out_valid(PE_8_io_data_0_out_valid),
    .io_data_0_out_bits(PE_8_io_data_0_out_bits)
  );
  PE PE_9 ( // @[pe.scala 184:13]
    .clock(PE_9_clock),
    .reset(PE_9_reset),
    .io_data_2_in_valid(PE_9_io_data_2_in_valid),
    .io_data_2_in_bits(PE_9_io_data_2_in_bits),
    .io_data_2_out_valid(PE_9_io_data_2_out_valid),
    .io_data_2_out_bits(PE_9_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_9_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_9_io_data_2_in_ready),
    .io_data_2_out_ready(PE_9_io_data_2_out_ready),
    .io_data_1_in_valid(PE_9_io_data_1_in_valid),
    .io_data_1_in_bits(PE_9_io_data_1_in_bits),
    .io_data_1_out_valid(PE_9_io_data_1_out_valid),
    .io_data_1_out_bits(PE_9_io_data_1_out_bits),
    .io_data_0_in_valid(PE_9_io_data_0_in_valid),
    .io_data_0_in_bits(PE_9_io_data_0_in_bits),
    .io_data_0_out_valid(PE_9_io_data_0_out_valid),
    .io_data_0_out_bits(PE_9_io_data_0_out_bits)
  );
  PE PE_10 ( // @[pe.scala 184:13]
    .clock(PE_10_clock),
    .reset(PE_10_reset),
    .io_data_2_in_valid(PE_10_io_data_2_in_valid),
    .io_data_2_in_bits(PE_10_io_data_2_in_bits),
    .io_data_2_out_valid(PE_10_io_data_2_out_valid),
    .io_data_2_out_bits(PE_10_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_10_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_10_io_data_2_in_ready),
    .io_data_2_out_ready(PE_10_io_data_2_out_ready),
    .io_data_1_in_valid(PE_10_io_data_1_in_valid),
    .io_data_1_in_bits(PE_10_io_data_1_in_bits),
    .io_data_1_out_valid(PE_10_io_data_1_out_valid),
    .io_data_1_out_bits(PE_10_io_data_1_out_bits),
    .io_data_0_in_valid(PE_10_io_data_0_in_valid),
    .io_data_0_in_bits(PE_10_io_data_0_in_bits),
    .io_data_0_out_valid(PE_10_io_data_0_out_valid),
    .io_data_0_out_bits(PE_10_io_data_0_out_bits)
  );
  PE PE_11 ( // @[pe.scala 184:13]
    .clock(PE_11_clock),
    .reset(PE_11_reset),
    .io_data_2_in_valid(PE_11_io_data_2_in_valid),
    .io_data_2_in_bits(PE_11_io_data_2_in_bits),
    .io_data_2_out_valid(PE_11_io_data_2_out_valid),
    .io_data_2_out_bits(PE_11_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_11_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_11_io_data_2_in_ready),
    .io_data_2_out_ready(PE_11_io_data_2_out_ready),
    .io_data_1_in_valid(PE_11_io_data_1_in_valid),
    .io_data_1_in_bits(PE_11_io_data_1_in_bits),
    .io_data_1_out_valid(PE_11_io_data_1_out_valid),
    .io_data_1_out_bits(PE_11_io_data_1_out_bits),
    .io_data_0_in_valid(PE_11_io_data_0_in_valid),
    .io_data_0_in_bits(PE_11_io_data_0_in_bits),
    .io_data_0_out_valid(PE_11_io_data_0_out_valid),
    .io_data_0_out_bits(PE_11_io_data_0_out_bits)
  );
  PE PE_12 ( // @[pe.scala 184:13]
    .clock(PE_12_clock),
    .reset(PE_12_reset),
    .io_data_2_in_valid(PE_12_io_data_2_in_valid),
    .io_data_2_in_bits(PE_12_io_data_2_in_bits),
    .io_data_2_out_valid(PE_12_io_data_2_out_valid),
    .io_data_2_out_bits(PE_12_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_12_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_12_io_data_2_in_ready),
    .io_data_2_out_ready(PE_12_io_data_2_out_ready),
    .io_data_1_in_valid(PE_12_io_data_1_in_valid),
    .io_data_1_in_bits(PE_12_io_data_1_in_bits),
    .io_data_1_out_valid(PE_12_io_data_1_out_valid),
    .io_data_1_out_bits(PE_12_io_data_1_out_bits),
    .io_data_0_in_valid(PE_12_io_data_0_in_valid),
    .io_data_0_in_bits(PE_12_io_data_0_in_bits),
    .io_data_0_out_valid(PE_12_io_data_0_out_valid),
    .io_data_0_out_bits(PE_12_io_data_0_out_bits)
  );
  PE PE_13 ( // @[pe.scala 184:13]
    .clock(PE_13_clock),
    .reset(PE_13_reset),
    .io_data_2_in_valid(PE_13_io_data_2_in_valid),
    .io_data_2_in_bits(PE_13_io_data_2_in_bits),
    .io_data_2_out_valid(PE_13_io_data_2_out_valid),
    .io_data_2_out_bits(PE_13_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_13_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_13_io_data_2_in_ready),
    .io_data_2_out_ready(PE_13_io_data_2_out_ready),
    .io_data_1_in_valid(PE_13_io_data_1_in_valid),
    .io_data_1_in_bits(PE_13_io_data_1_in_bits),
    .io_data_1_out_valid(PE_13_io_data_1_out_valid),
    .io_data_1_out_bits(PE_13_io_data_1_out_bits),
    .io_data_0_in_valid(PE_13_io_data_0_in_valid),
    .io_data_0_in_bits(PE_13_io_data_0_in_bits),
    .io_data_0_out_valid(PE_13_io_data_0_out_valid),
    .io_data_0_out_bits(PE_13_io_data_0_out_bits)
  );
  PE PE_14 ( // @[pe.scala 184:13]
    .clock(PE_14_clock),
    .reset(PE_14_reset),
    .io_data_2_in_valid(PE_14_io_data_2_in_valid),
    .io_data_2_in_bits(PE_14_io_data_2_in_bits),
    .io_data_2_out_valid(PE_14_io_data_2_out_valid),
    .io_data_2_out_bits(PE_14_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_14_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_14_io_data_2_in_ready),
    .io_data_2_out_ready(PE_14_io_data_2_out_ready),
    .io_data_1_in_valid(PE_14_io_data_1_in_valid),
    .io_data_1_in_bits(PE_14_io_data_1_in_bits),
    .io_data_1_out_valid(PE_14_io_data_1_out_valid),
    .io_data_1_out_bits(PE_14_io_data_1_out_bits),
    .io_data_0_in_valid(PE_14_io_data_0_in_valid),
    .io_data_0_in_bits(PE_14_io_data_0_in_bits),
    .io_data_0_out_valid(PE_14_io_data_0_out_valid),
    .io_data_0_out_bits(PE_14_io_data_0_out_bits)
  );
  PE PE_15 ( // @[pe.scala 184:13]
    .clock(PE_15_clock),
    .reset(PE_15_reset),
    .io_data_2_in_valid(PE_15_io_data_2_in_valid),
    .io_data_2_in_bits(PE_15_io_data_2_in_bits),
    .io_data_2_out_valid(PE_15_io_data_2_out_valid),
    .io_data_2_out_bits(PE_15_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_15_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_15_io_data_2_in_ready),
    .io_data_2_out_ready(PE_15_io_data_2_out_ready),
    .io_data_1_in_valid(PE_15_io_data_1_in_valid),
    .io_data_1_in_bits(PE_15_io_data_1_in_bits),
    .io_data_1_out_valid(PE_15_io_data_1_out_valid),
    .io_data_1_out_bits(PE_15_io_data_1_out_bits),
    .io_data_0_in_valid(PE_15_io_data_0_in_valid),
    .io_data_0_in_bits(PE_15_io_data_0_in_bits),
    .io_data_0_out_valid(PE_15_io_data_0_out_valid),
    .io_data_0_out_bits(PE_15_io_data_0_out_bits)
  );
  PE PE_16 ( // @[pe.scala 184:13]
    .clock(PE_16_clock),
    .reset(PE_16_reset),
    .io_data_2_in_valid(PE_16_io_data_2_in_valid),
    .io_data_2_in_bits(PE_16_io_data_2_in_bits),
    .io_data_2_out_valid(PE_16_io_data_2_out_valid),
    .io_data_2_out_bits(PE_16_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_16_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_16_io_data_2_in_ready),
    .io_data_2_out_ready(PE_16_io_data_2_out_ready),
    .io_data_1_in_valid(PE_16_io_data_1_in_valid),
    .io_data_1_in_bits(PE_16_io_data_1_in_bits),
    .io_data_1_out_valid(PE_16_io_data_1_out_valid),
    .io_data_1_out_bits(PE_16_io_data_1_out_bits),
    .io_data_0_in_valid(PE_16_io_data_0_in_valid),
    .io_data_0_in_bits(PE_16_io_data_0_in_bits),
    .io_data_0_out_valid(PE_16_io_data_0_out_valid),
    .io_data_0_out_bits(PE_16_io_data_0_out_bits)
  );
  PE PE_17 ( // @[pe.scala 184:13]
    .clock(PE_17_clock),
    .reset(PE_17_reset),
    .io_data_2_in_valid(PE_17_io_data_2_in_valid),
    .io_data_2_in_bits(PE_17_io_data_2_in_bits),
    .io_data_2_out_valid(PE_17_io_data_2_out_valid),
    .io_data_2_out_bits(PE_17_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_17_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_17_io_data_2_in_ready),
    .io_data_2_out_ready(PE_17_io_data_2_out_ready),
    .io_data_1_in_valid(PE_17_io_data_1_in_valid),
    .io_data_1_in_bits(PE_17_io_data_1_in_bits),
    .io_data_1_out_valid(PE_17_io_data_1_out_valid),
    .io_data_1_out_bits(PE_17_io_data_1_out_bits),
    .io_data_0_in_valid(PE_17_io_data_0_in_valid),
    .io_data_0_in_bits(PE_17_io_data_0_in_bits),
    .io_data_0_out_valid(PE_17_io_data_0_out_valid),
    .io_data_0_out_bits(PE_17_io_data_0_out_bits)
  );
  PE PE_18 ( // @[pe.scala 184:13]
    .clock(PE_18_clock),
    .reset(PE_18_reset),
    .io_data_2_in_valid(PE_18_io_data_2_in_valid),
    .io_data_2_in_bits(PE_18_io_data_2_in_bits),
    .io_data_2_out_valid(PE_18_io_data_2_out_valid),
    .io_data_2_out_bits(PE_18_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_18_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_18_io_data_2_in_ready),
    .io_data_2_out_ready(PE_18_io_data_2_out_ready),
    .io_data_1_in_valid(PE_18_io_data_1_in_valid),
    .io_data_1_in_bits(PE_18_io_data_1_in_bits),
    .io_data_1_out_valid(PE_18_io_data_1_out_valid),
    .io_data_1_out_bits(PE_18_io_data_1_out_bits),
    .io_data_0_in_valid(PE_18_io_data_0_in_valid),
    .io_data_0_in_bits(PE_18_io_data_0_in_bits),
    .io_data_0_out_valid(PE_18_io_data_0_out_valid),
    .io_data_0_out_bits(PE_18_io_data_0_out_bits)
  );
  PE PE_19 ( // @[pe.scala 184:13]
    .clock(PE_19_clock),
    .reset(PE_19_reset),
    .io_data_2_in_valid(PE_19_io_data_2_in_valid),
    .io_data_2_in_bits(PE_19_io_data_2_in_bits),
    .io_data_2_out_valid(PE_19_io_data_2_out_valid),
    .io_data_2_out_bits(PE_19_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_19_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_19_io_data_2_in_ready),
    .io_data_2_out_ready(PE_19_io_data_2_out_ready),
    .io_data_1_in_valid(PE_19_io_data_1_in_valid),
    .io_data_1_in_bits(PE_19_io_data_1_in_bits),
    .io_data_1_out_valid(PE_19_io_data_1_out_valid),
    .io_data_1_out_bits(PE_19_io_data_1_out_bits),
    .io_data_0_in_valid(PE_19_io_data_0_in_valid),
    .io_data_0_in_bits(PE_19_io_data_0_in_bits),
    .io_data_0_out_valid(PE_19_io_data_0_out_valid),
    .io_data_0_out_bits(PE_19_io_data_0_out_bits)
  );
  PE PE_20 ( // @[pe.scala 184:13]
    .clock(PE_20_clock),
    .reset(PE_20_reset),
    .io_data_2_in_valid(PE_20_io_data_2_in_valid),
    .io_data_2_in_bits(PE_20_io_data_2_in_bits),
    .io_data_2_out_valid(PE_20_io_data_2_out_valid),
    .io_data_2_out_bits(PE_20_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_20_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_20_io_data_2_in_ready),
    .io_data_2_out_ready(PE_20_io_data_2_out_ready),
    .io_data_1_in_valid(PE_20_io_data_1_in_valid),
    .io_data_1_in_bits(PE_20_io_data_1_in_bits),
    .io_data_1_out_valid(PE_20_io_data_1_out_valid),
    .io_data_1_out_bits(PE_20_io_data_1_out_bits),
    .io_data_0_in_valid(PE_20_io_data_0_in_valid),
    .io_data_0_in_bits(PE_20_io_data_0_in_bits),
    .io_data_0_out_valid(PE_20_io_data_0_out_valid),
    .io_data_0_out_bits(PE_20_io_data_0_out_bits)
  );
  PE PE_21 ( // @[pe.scala 184:13]
    .clock(PE_21_clock),
    .reset(PE_21_reset),
    .io_data_2_in_valid(PE_21_io_data_2_in_valid),
    .io_data_2_in_bits(PE_21_io_data_2_in_bits),
    .io_data_2_out_valid(PE_21_io_data_2_out_valid),
    .io_data_2_out_bits(PE_21_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_21_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_21_io_data_2_in_ready),
    .io_data_2_out_ready(PE_21_io_data_2_out_ready),
    .io_data_1_in_valid(PE_21_io_data_1_in_valid),
    .io_data_1_in_bits(PE_21_io_data_1_in_bits),
    .io_data_1_out_valid(PE_21_io_data_1_out_valid),
    .io_data_1_out_bits(PE_21_io_data_1_out_bits),
    .io_data_0_in_valid(PE_21_io_data_0_in_valid),
    .io_data_0_in_bits(PE_21_io_data_0_in_bits),
    .io_data_0_out_valid(PE_21_io_data_0_out_valid),
    .io_data_0_out_bits(PE_21_io_data_0_out_bits)
  );
  PE PE_22 ( // @[pe.scala 184:13]
    .clock(PE_22_clock),
    .reset(PE_22_reset),
    .io_data_2_in_valid(PE_22_io_data_2_in_valid),
    .io_data_2_in_bits(PE_22_io_data_2_in_bits),
    .io_data_2_out_valid(PE_22_io_data_2_out_valid),
    .io_data_2_out_bits(PE_22_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_22_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_22_io_data_2_in_ready),
    .io_data_2_out_ready(PE_22_io_data_2_out_ready),
    .io_data_1_in_valid(PE_22_io_data_1_in_valid),
    .io_data_1_in_bits(PE_22_io_data_1_in_bits),
    .io_data_1_out_valid(PE_22_io_data_1_out_valid),
    .io_data_1_out_bits(PE_22_io_data_1_out_bits),
    .io_data_0_in_valid(PE_22_io_data_0_in_valid),
    .io_data_0_in_bits(PE_22_io_data_0_in_bits),
    .io_data_0_out_valid(PE_22_io_data_0_out_valid),
    .io_data_0_out_bits(PE_22_io_data_0_out_bits)
  );
  PE PE_23 ( // @[pe.scala 184:13]
    .clock(PE_23_clock),
    .reset(PE_23_reset),
    .io_data_2_in_valid(PE_23_io_data_2_in_valid),
    .io_data_2_in_bits(PE_23_io_data_2_in_bits),
    .io_data_2_out_valid(PE_23_io_data_2_out_valid),
    .io_data_2_out_bits(PE_23_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_23_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_23_io_data_2_in_ready),
    .io_data_2_out_ready(PE_23_io_data_2_out_ready),
    .io_data_1_in_valid(PE_23_io_data_1_in_valid),
    .io_data_1_in_bits(PE_23_io_data_1_in_bits),
    .io_data_1_out_valid(PE_23_io_data_1_out_valid),
    .io_data_1_out_bits(PE_23_io_data_1_out_bits),
    .io_data_0_in_valid(PE_23_io_data_0_in_valid),
    .io_data_0_in_bits(PE_23_io_data_0_in_bits),
    .io_data_0_out_valid(PE_23_io_data_0_out_valid),
    .io_data_0_out_bits(PE_23_io_data_0_out_bits)
  );
  PE PE_24 ( // @[pe.scala 184:13]
    .clock(PE_24_clock),
    .reset(PE_24_reset),
    .io_data_2_in_valid(PE_24_io_data_2_in_valid),
    .io_data_2_in_bits(PE_24_io_data_2_in_bits),
    .io_data_2_out_valid(PE_24_io_data_2_out_valid),
    .io_data_2_out_bits(PE_24_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_24_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_24_io_data_2_in_ready),
    .io_data_2_out_ready(PE_24_io_data_2_out_ready),
    .io_data_1_in_valid(PE_24_io_data_1_in_valid),
    .io_data_1_in_bits(PE_24_io_data_1_in_bits),
    .io_data_1_out_valid(PE_24_io_data_1_out_valid),
    .io_data_1_out_bits(PE_24_io_data_1_out_bits),
    .io_data_0_in_valid(PE_24_io_data_0_in_valid),
    .io_data_0_in_bits(PE_24_io_data_0_in_bits),
    .io_data_0_out_valid(PE_24_io_data_0_out_valid),
    .io_data_0_out_bits(PE_24_io_data_0_out_bits)
  );
  PE PE_25 ( // @[pe.scala 184:13]
    .clock(PE_25_clock),
    .reset(PE_25_reset),
    .io_data_2_in_valid(PE_25_io_data_2_in_valid),
    .io_data_2_in_bits(PE_25_io_data_2_in_bits),
    .io_data_2_out_valid(PE_25_io_data_2_out_valid),
    .io_data_2_out_bits(PE_25_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_25_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_25_io_data_2_in_ready),
    .io_data_2_out_ready(PE_25_io_data_2_out_ready),
    .io_data_1_in_valid(PE_25_io_data_1_in_valid),
    .io_data_1_in_bits(PE_25_io_data_1_in_bits),
    .io_data_1_out_valid(PE_25_io_data_1_out_valid),
    .io_data_1_out_bits(PE_25_io_data_1_out_bits),
    .io_data_0_in_valid(PE_25_io_data_0_in_valid),
    .io_data_0_in_bits(PE_25_io_data_0_in_bits),
    .io_data_0_out_valid(PE_25_io_data_0_out_valid),
    .io_data_0_out_bits(PE_25_io_data_0_out_bits)
  );
  PE PE_26 ( // @[pe.scala 184:13]
    .clock(PE_26_clock),
    .reset(PE_26_reset),
    .io_data_2_in_valid(PE_26_io_data_2_in_valid),
    .io_data_2_in_bits(PE_26_io_data_2_in_bits),
    .io_data_2_out_valid(PE_26_io_data_2_out_valid),
    .io_data_2_out_bits(PE_26_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_26_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_26_io_data_2_in_ready),
    .io_data_2_out_ready(PE_26_io_data_2_out_ready),
    .io_data_1_in_valid(PE_26_io_data_1_in_valid),
    .io_data_1_in_bits(PE_26_io_data_1_in_bits),
    .io_data_1_out_valid(PE_26_io_data_1_out_valid),
    .io_data_1_out_bits(PE_26_io_data_1_out_bits),
    .io_data_0_in_valid(PE_26_io_data_0_in_valid),
    .io_data_0_in_bits(PE_26_io_data_0_in_bits),
    .io_data_0_out_valid(PE_26_io_data_0_out_valid),
    .io_data_0_out_bits(PE_26_io_data_0_out_bits)
  );
  PE PE_27 ( // @[pe.scala 184:13]
    .clock(PE_27_clock),
    .reset(PE_27_reset),
    .io_data_2_in_valid(PE_27_io_data_2_in_valid),
    .io_data_2_in_bits(PE_27_io_data_2_in_bits),
    .io_data_2_out_valid(PE_27_io_data_2_out_valid),
    .io_data_2_out_bits(PE_27_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_27_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_27_io_data_2_in_ready),
    .io_data_2_out_ready(PE_27_io_data_2_out_ready),
    .io_data_1_in_valid(PE_27_io_data_1_in_valid),
    .io_data_1_in_bits(PE_27_io_data_1_in_bits),
    .io_data_1_out_valid(PE_27_io_data_1_out_valid),
    .io_data_1_out_bits(PE_27_io_data_1_out_bits),
    .io_data_0_in_valid(PE_27_io_data_0_in_valid),
    .io_data_0_in_bits(PE_27_io_data_0_in_bits),
    .io_data_0_out_valid(PE_27_io_data_0_out_valid),
    .io_data_0_out_bits(PE_27_io_data_0_out_bits)
  );
  PE PE_28 ( // @[pe.scala 184:13]
    .clock(PE_28_clock),
    .reset(PE_28_reset),
    .io_data_2_in_valid(PE_28_io_data_2_in_valid),
    .io_data_2_in_bits(PE_28_io_data_2_in_bits),
    .io_data_2_out_valid(PE_28_io_data_2_out_valid),
    .io_data_2_out_bits(PE_28_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_28_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_28_io_data_2_in_ready),
    .io_data_2_out_ready(PE_28_io_data_2_out_ready),
    .io_data_1_in_valid(PE_28_io_data_1_in_valid),
    .io_data_1_in_bits(PE_28_io_data_1_in_bits),
    .io_data_1_out_valid(PE_28_io_data_1_out_valid),
    .io_data_1_out_bits(PE_28_io_data_1_out_bits),
    .io_data_0_in_valid(PE_28_io_data_0_in_valid),
    .io_data_0_in_bits(PE_28_io_data_0_in_bits),
    .io_data_0_out_valid(PE_28_io_data_0_out_valid),
    .io_data_0_out_bits(PE_28_io_data_0_out_bits)
  );
  PE PE_29 ( // @[pe.scala 184:13]
    .clock(PE_29_clock),
    .reset(PE_29_reset),
    .io_data_2_in_valid(PE_29_io_data_2_in_valid),
    .io_data_2_in_bits(PE_29_io_data_2_in_bits),
    .io_data_2_out_valid(PE_29_io_data_2_out_valid),
    .io_data_2_out_bits(PE_29_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_29_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_29_io_data_2_in_ready),
    .io_data_2_out_ready(PE_29_io_data_2_out_ready),
    .io_data_1_in_valid(PE_29_io_data_1_in_valid),
    .io_data_1_in_bits(PE_29_io_data_1_in_bits),
    .io_data_1_out_valid(PE_29_io_data_1_out_valid),
    .io_data_1_out_bits(PE_29_io_data_1_out_bits),
    .io_data_0_in_valid(PE_29_io_data_0_in_valid),
    .io_data_0_in_bits(PE_29_io_data_0_in_bits),
    .io_data_0_out_valid(PE_29_io_data_0_out_valid),
    .io_data_0_out_bits(PE_29_io_data_0_out_bits)
  );
  PE PE_30 ( // @[pe.scala 184:13]
    .clock(PE_30_clock),
    .reset(PE_30_reset),
    .io_data_2_in_valid(PE_30_io_data_2_in_valid),
    .io_data_2_in_bits(PE_30_io_data_2_in_bits),
    .io_data_2_out_valid(PE_30_io_data_2_out_valid),
    .io_data_2_out_bits(PE_30_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_30_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_30_io_data_2_in_ready),
    .io_data_2_out_ready(PE_30_io_data_2_out_ready),
    .io_data_1_in_valid(PE_30_io_data_1_in_valid),
    .io_data_1_in_bits(PE_30_io_data_1_in_bits),
    .io_data_1_out_valid(PE_30_io_data_1_out_valid),
    .io_data_1_out_bits(PE_30_io_data_1_out_bits),
    .io_data_0_in_valid(PE_30_io_data_0_in_valid),
    .io_data_0_in_bits(PE_30_io_data_0_in_bits),
    .io_data_0_out_valid(PE_30_io_data_0_out_valid),
    .io_data_0_out_bits(PE_30_io_data_0_out_bits)
  );
  PE PE_31 ( // @[pe.scala 184:13]
    .clock(PE_31_clock),
    .reset(PE_31_reset),
    .io_data_2_in_valid(PE_31_io_data_2_in_valid),
    .io_data_2_in_bits(PE_31_io_data_2_in_bits),
    .io_data_2_out_valid(PE_31_io_data_2_out_valid),
    .io_data_2_out_bits(PE_31_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_31_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_31_io_data_2_in_ready),
    .io_data_2_out_ready(PE_31_io_data_2_out_ready),
    .io_data_1_in_valid(PE_31_io_data_1_in_valid),
    .io_data_1_in_bits(PE_31_io_data_1_in_bits),
    .io_data_1_out_valid(PE_31_io_data_1_out_valid),
    .io_data_1_out_bits(PE_31_io_data_1_out_bits),
    .io_data_0_in_valid(PE_31_io_data_0_in_valid),
    .io_data_0_in_bits(PE_31_io_data_0_in_bits),
    .io_data_0_out_valid(PE_31_io_data_0_out_valid),
    .io_data_0_out_bits(PE_31_io_data_0_out_bits)
  );
  PE PE_32 ( // @[pe.scala 184:13]
    .clock(PE_32_clock),
    .reset(PE_32_reset),
    .io_data_2_in_valid(PE_32_io_data_2_in_valid),
    .io_data_2_in_bits(PE_32_io_data_2_in_bits),
    .io_data_2_out_valid(PE_32_io_data_2_out_valid),
    .io_data_2_out_bits(PE_32_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_32_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_32_io_data_2_in_ready),
    .io_data_2_out_ready(PE_32_io_data_2_out_ready),
    .io_data_1_in_valid(PE_32_io_data_1_in_valid),
    .io_data_1_in_bits(PE_32_io_data_1_in_bits),
    .io_data_1_out_valid(PE_32_io_data_1_out_valid),
    .io_data_1_out_bits(PE_32_io_data_1_out_bits),
    .io_data_0_in_valid(PE_32_io_data_0_in_valid),
    .io_data_0_in_bits(PE_32_io_data_0_in_bits),
    .io_data_0_out_valid(PE_32_io_data_0_out_valid),
    .io_data_0_out_bits(PE_32_io_data_0_out_bits)
  );
  PE PE_33 ( // @[pe.scala 184:13]
    .clock(PE_33_clock),
    .reset(PE_33_reset),
    .io_data_2_in_valid(PE_33_io_data_2_in_valid),
    .io_data_2_in_bits(PE_33_io_data_2_in_bits),
    .io_data_2_out_valid(PE_33_io_data_2_out_valid),
    .io_data_2_out_bits(PE_33_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_33_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_33_io_data_2_in_ready),
    .io_data_2_out_ready(PE_33_io_data_2_out_ready),
    .io_data_1_in_valid(PE_33_io_data_1_in_valid),
    .io_data_1_in_bits(PE_33_io_data_1_in_bits),
    .io_data_1_out_valid(PE_33_io_data_1_out_valid),
    .io_data_1_out_bits(PE_33_io_data_1_out_bits),
    .io_data_0_in_valid(PE_33_io_data_0_in_valid),
    .io_data_0_in_bits(PE_33_io_data_0_in_bits),
    .io_data_0_out_valid(PE_33_io_data_0_out_valid),
    .io_data_0_out_bits(PE_33_io_data_0_out_bits)
  );
  PE PE_34 ( // @[pe.scala 184:13]
    .clock(PE_34_clock),
    .reset(PE_34_reset),
    .io_data_2_in_valid(PE_34_io_data_2_in_valid),
    .io_data_2_in_bits(PE_34_io_data_2_in_bits),
    .io_data_2_out_valid(PE_34_io_data_2_out_valid),
    .io_data_2_out_bits(PE_34_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_34_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_34_io_data_2_in_ready),
    .io_data_2_out_ready(PE_34_io_data_2_out_ready),
    .io_data_1_in_valid(PE_34_io_data_1_in_valid),
    .io_data_1_in_bits(PE_34_io_data_1_in_bits),
    .io_data_1_out_valid(PE_34_io_data_1_out_valid),
    .io_data_1_out_bits(PE_34_io_data_1_out_bits),
    .io_data_0_in_valid(PE_34_io_data_0_in_valid),
    .io_data_0_in_bits(PE_34_io_data_0_in_bits),
    .io_data_0_out_valid(PE_34_io_data_0_out_valid),
    .io_data_0_out_bits(PE_34_io_data_0_out_bits)
  );
  PE PE_35 ( // @[pe.scala 184:13]
    .clock(PE_35_clock),
    .reset(PE_35_reset),
    .io_data_2_in_valid(PE_35_io_data_2_in_valid),
    .io_data_2_in_bits(PE_35_io_data_2_in_bits),
    .io_data_2_out_valid(PE_35_io_data_2_out_valid),
    .io_data_2_out_bits(PE_35_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_35_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_35_io_data_2_in_ready),
    .io_data_2_out_ready(PE_35_io_data_2_out_ready),
    .io_data_1_in_valid(PE_35_io_data_1_in_valid),
    .io_data_1_in_bits(PE_35_io_data_1_in_bits),
    .io_data_1_out_valid(PE_35_io_data_1_out_valid),
    .io_data_1_out_bits(PE_35_io_data_1_out_bits),
    .io_data_0_in_valid(PE_35_io_data_0_in_valid),
    .io_data_0_in_bits(PE_35_io_data_0_in_bits),
    .io_data_0_out_valid(PE_35_io_data_0_out_valid),
    .io_data_0_out_bits(PE_35_io_data_0_out_bits)
  );
  PE PE_36 ( // @[pe.scala 184:13]
    .clock(PE_36_clock),
    .reset(PE_36_reset),
    .io_data_2_in_valid(PE_36_io_data_2_in_valid),
    .io_data_2_in_bits(PE_36_io_data_2_in_bits),
    .io_data_2_out_valid(PE_36_io_data_2_out_valid),
    .io_data_2_out_bits(PE_36_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_36_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_36_io_data_2_in_ready),
    .io_data_2_out_ready(PE_36_io_data_2_out_ready),
    .io_data_1_in_valid(PE_36_io_data_1_in_valid),
    .io_data_1_in_bits(PE_36_io_data_1_in_bits),
    .io_data_1_out_valid(PE_36_io_data_1_out_valid),
    .io_data_1_out_bits(PE_36_io_data_1_out_bits),
    .io_data_0_in_valid(PE_36_io_data_0_in_valid),
    .io_data_0_in_bits(PE_36_io_data_0_in_bits),
    .io_data_0_out_valid(PE_36_io_data_0_out_valid),
    .io_data_0_out_bits(PE_36_io_data_0_out_bits)
  );
  PE PE_37 ( // @[pe.scala 184:13]
    .clock(PE_37_clock),
    .reset(PE_37_reset),
    .io_data_2_in_valid(PE_37_io_data_2_in_valid),
    .io_data_2_in_bits(PE_37_io_data_2_in_bits),
    .io_data_2_out_valid(PE_37_io_data_2_out_valid),
    .io_data_2_out_bits(PE_37_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_37_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_37_io_data_2_in_ready),
    .io_data_2_out_ready(PE_37_io_data_2_out_ready),
    .io_data_1_in_valid(PE_37_io_data_1_in_valid),
    .io_data_1_in_bits(PE_37_io_data_1_in_bits),
    .io_data_1_out_valid(PE_37_io_data_1_out_valid),
    .io_data_1_out_bits(PE_37_io_data_1_out_bits),
    .io_data_0_in_valid(PE_37_io_data_0_in_valid),
    .io_data_0_in_bits(PE_37_io_data_0_in_bits),
    .io_data_0_out_valid(PE_37_io_data_0_out_valid),
    .io_data_0_out_bits(PE_37_io_data_0_out_bits)
  );
  PE PE_38 ( // @[pe.scala 184:13]
    .clock(PE_38_clock),
    .reset(PE_38_reset),
    .io_data_2_in_valid(PE_38_io_data_2_in_valid),
    .io_data_2_in_bits(PE_38_io_data_2_in_bits),
    .io_data_2_out_valid(PE_38_io_data_2_out_valid),
    .io_data_2_out_bits(PE_38_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_38_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_38_io_data_2_in_ready),
    .io_data_2_out_ready(PE_38_io_data_2_out_ready),
    .io_data_1_in_valid(PE_38_io_data_1_in_valid),
    .io_data_1_in_bits(PE_38_io_data_1_in_bits),
    .io_data_1_out_valid(PE_38_io_data_1_out_valid),
    .io_data_1_out_bits(PE_38_io_data_1_out_bits),
    .io_data_0_in_valid(PE_38_io_data_0_in_valid),
    .io_data_0_in_bits(PE_38_io_data_0_in_bits),
    .io_data_0_out_valid(PE_38_io_data_0_out_valid),
    .io_data_0_out_bits(PE_38_io_data_0_out_bits)
  );
  PE PE_39 ( // @[pe.scala 184:13]
    .clock(PE_39_clock),
    .reset(PE_39_reset),
    .io_data_2_in_valid(PE_39_io_data_2_in_valid),
    .io_data_2_in_bits(PE_39_io_data_2_in_bits),
    .io_data_2_out_valid(PE_39_io_data_2_out_valid),
    .io_data_2_out_bits(PE_39_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_39_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_39_io_data_2_in_ready),
    .io_data_2_out_ready(PE_39_io_data_2_out_ready),
    .io_data_1_in_valid(PE_39_io_data_1_in_valid),
    .io_data_1_in_bits(PE_39_io_data_1_in_bits),
    .io_data_1_out_valid(PE_39_io_data_1_out_valid),
    .io_data_1_out_bits(PE_39_io_data_1_out_bits),
    .io_data_0_in_valid(PE_39_io_data_0_in_valid),
    .io_data_0_in_bits(PE_39_io_data_0_in_bits),
    .io_data_0_out_valid(PE_39_io_data_0_out_valid),
    .io_data_0_out_bits(PE_39_io_data_0_out_bits)
  );
  PE PE_40 ( // @[pe.scala 184:13]
    .clock(PE_40_clock),
    .reset(PE_40_reset),
    .io_data_2_in_valid(PE_40_io_data_2_in_valid),
    .io_data_2_in_bits(PE_40_io_data_2_in_bits),
    .io_data_2_out_valid(PE_40_io_data_2_out_valid),
    .io_data_2_out_bits(PE_40_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_40_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_40_io_data_2_in_ready),
    .io_data_2_out_ready(PE_40_io_data_2_out_ready),
    .io_data_1_in_valid(PE_40_io_data_1_in_valid),
    .io_data_1_in_bits(PE_40_io_data_1_in_bits),
    .io_data_1_out_valid(PE_40_io_data_1_out_valid),
    .io_data_1_out_bits(PE_40_io_data_1_out_bits),
    .io_data_0_in_valid(PE_40_io_data_0_in_valid),
    .io_data_0_in_bits(PE_40_io_data_0_in_bits),
    .io_data_0_out_valid(PE_40_io_data_0_out_valid),
    .io_data_0_out_bits(PE_40_io_data_0_out_bits)
  );
  PE PE_41 ( // @[pe.scala 184:13]
    .clock(PE_41_clock),
    .reset(PE_41_reset),
    .io_data_2_in_valid(PE_41_io_data_2_in_valid),
    .io_data_2_in_bits(PE_41_io_data_2_in_bits),
    .io_data_2_out_valid(PE_41_io_data_2_out_valid),
    .io_data_2_out_bits(PE_41_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_41_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_41_io_data_2_in_ready),
    .io_data_2_out_ready(PE_41_io_data_2_out_ready),
    .io_data_1_in_valid(PE_41_io_data_1_in_valid),
    .io_data_1_in_bits(PE_41_io_data_1_in_bits),
    .io_data_1_out_valid(PE_41_io_data_1_out_valid),
    .io_data_1_out_bits(PE_41_io_data_1_out_bits),
    .io_data_0_in_valid(PE_41_io_data_0_in_valid),
    .io_data_0_in_bits(PE_41_io_data_0_in_bits),
    .io_data_0_out_valid(PE_41_io_data_0_out_valid),
    .io_data_0_out_bits(PE_41_io_data_0_out_bits)
  );
  PE PE_42 ( // @[pe.scala 184:13]
    .clock(PE_42_clock),
    .reset(PE_42_reset),
    .io_data_2_in_valid(PE_42_io_data_2_in_valid),
    .io_data_2_in_bits(PE_42_io_data_2_in_bits),
    .io_data_2_out_valid(PE_42_io_data_2_out_valid),
    .io_data_2_out_bits(PE_42_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_42_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_42_io_data_2_in_ready),
    .io_data_2_out_ready(PE_42_io_data_2_out_ready),
    .io_data_1_in_valid(PE_42_io_data_1_in_valid),
    .io_data_1_in_bits(PE_42_io_data_1_in_bits),
    .io_data_1_out_valid(PE_42_io_data_1_out_valid),
    .io_data_1_out_bits(PE_42_io_data_1_out_bits),
    .io_data_0_in_valid(PE_42_io_data_0_in_valid),
    .io_data_0_in_bits(PE_42_io_data_0_in_bits),
    .io_data_0_out_valid(PE_42_io_data_0_out_valid),
    .io_data_0_out_bits(PE_42_io_data_0_out_bits)
  );
  PE PE_43 ( // @[pe.scala 184:13]
    .clock(PE_43_clock),
    .reset(PE_43_reset),
    .io_data_2_in_valid(PE_43_io_data_2_in_valid),
    .io_data_2_in_bits(PE_43_io_data_2_in_bits),
    .io_data_2_out_valid(PE_43_io_data_2_out_valid),
    .io_data_2_out_bits(PE_43_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_43_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_43_io_data_2_in_ready),
    .io_data_2_out_ready(PE_43_io_data_2_out_ready),
    .io_data_1_in_valid(PE_43_io_data_1_in_valid),
    .io_data_1_in_bits(PE_43_io_data_1_in_bits),
    .io_data_1_out_valid(PE_43_io_data_1_out_valid),
    .io_data_1_out_bits(PE_43_io_data_1_out_bits),
    .io_data_0_in_valid(PE_43_io_data_0_in_valid),
    .io_data_0_in_bits(PE_43_io_data_0_in_bits),
    .io_data_0_out_valid(PE_43_io_data_0_out_valid),
    .io_data_0_out_bits(PE_43_io_data_0_out_bits)
  );
  PE PE_44 ( // @[pe.scala 184:13]
    .clock(PE_44_clock),
    .reset(PE_44_reset),
    .io_data_2_in_valid(PE_44_io_data_2_in_valid),
    .io_data_2_in_bits(PE_44_io_data_2_in_bits),
    .io_data_2_out_valid(PE_44_io_data_2_out_valid),
    .io_data_2_out_bits(PE_44_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_44_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_44_io_data_2_in_ready),
    .io_data_2_out_ready(PE_44_io_data_2_out_ready),
    .io_data_1_in_valid(PE_44_io_data_1_in_valid),
    .io_data_1_in_bits(PE_44_io_data_1_in_bits),
    .io_data_1_out_valid(PE_44_io_data_1_out_valid),
    .io_data_1_out_bits(PE_44_io_data_1_out_bits),
    .io_data_0_in_valid(PE_44_io_data_0_in_valid),
    .io_data_0_in_bits(PE_44_io_data_0_in_bits),
    .io_data_0_out_valid(PE_44_io_data_0_out_valid),
    .io_data_0_out_bits(PE_44_io_data_0_out_bits)
  );
  PE PE_45 ( // @[pe.scala 184:13]
    .clock(PE_45_clock),
    .reset(PE_45_reset),
    .io_data_2_in_valid(PE_45_io_data_2_in_valid),
    .io_data_2_in_bits(PE_45_io_data_2_in_bits),
    .io_data_2_out_valid(PE_45_io_data_2_out_valid),
    .io_data_2_out_bits(PE_45_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_45_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_45_io_data_2_in_ready),
    .io_data_2_out_ready(PE_45_io_data_2_out_ready),
    .io_data_1_in_valid(PE_45_io_data_1_in_valid),
    .io_data_1_in_bits(PE_45_io_data_1_in_bits),
    .io_data_1_out_valid(PE_45_io_data_1_out_valid),
    .io_data_1_out_bits(PE_45_io_data_1_out_bits),
    .io_data_0_in_valid(PE_45_io_data_0_in_valid),
    .io_data_0_in_bits(PE_45_io_data_0_in_bits),
    .io_data_0_out_valid(PE_45_io_data_0_out_valid),
    .io_data_0_out_bits(PE_45_io_data_0_out_bits)
  );
  PE PE_46 ( // @[pe.scala 184:13]
    .clock(PE_46_clock),
    .reset(PE_46_reset),
    .io_data_2_in_valid(PE_46_io_data_2_in_valid),
    .io_data_2_in_bits(PE_46_io_data_2_in_bits),
    .io_data_2_out_valid(PE_46_io_data_2_out_valid),
    .io_data_2_out_bits(PE_46_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_46_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_46_io_data_2_in_ready),
    .io_data_2_out_ready(PE_46_io_data_2_out_ready),
    .io_data_1_in_valid(PE_46_io_data_1_in_valid),
    .io_data_1_in_bits(PE_46_io_data_1_in_bits),
    .io_data_1_out_valid(PE_46_io_data_1_out_valid),
    .io_data_1_out_bits(PE_46_io_data_1_out_bits),
    .io_data_0_in_valid(PE_46_io_data_0_in_valid),
    .io_data_0_in_bits(PE_46_io_data_0_in_bits),
    .io_data_0_out_valid(PE_46_io_data_0_out_valid),
    .io_data_0_out_bits(PE_46_io_data_0_out_bits)
  );
  PE PE_47 ( // @[pe.scala 184:13]
    .clock(PE_47_clock),
    .reset(PE_47_reset),
    .io_data_2_in_valid(PE_47_io_data_2_in_valid),
    .io_data_2_in_bits(PE_47_io_data_2_in_bits),
    .io_data_2_out_valid(PE_47_io_data_2_out_valid),
    .io_data_2_out_bits(PE_47_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_47_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_47_io_data_2_in_ready),
    .io_data_2_out_ready(PE_47_io_data_2_out_ready),
    .io_data_1_in_valid(PE_47_io_data_1_in_valid),
    .io_data_1_in_bits(PE_47_io_data_1_in_bits),
    .io_data_1_out_valid(PE_47_io_data_1_out_valid),
    .io_data_1_out_bits(PE_47_io_data_1_out_bits),
    .io_data_0_in_valid(PE_47_io_data_0_in_valid),
    .io_data_0_in_bits(PE_47_io_data_0_in_bits),
    .io_data_0_out_valid(PE_47_io_data_0_out_valid),
    .io_data_0_out_bits(PE_47_io_data_0_out_bits)
  );
  PE PE_48 ( // @[pe.scala 184:13]
    .clock(PE_48_clock),
    .reset(PE_48_reset),
    .io_data_2_in_valid(PE_48_io_data_2_in_valid),
    .io_data_2_in_bits(PE_48_io_data_2_in_bits),
    .io_data_2_out_valid(PE_48_io_data_2_out_valid),
    .io_data_2_out_bits(PE_48_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_48_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_48_io_data_2_in_ready),
    .io_data_2_out_ready(PE_48_io_data_2_out_ready),
    .io_data_1_in_valid(PE_48_io_data_1_in_valid),
    .io_data_1_in_bits(PE_48_io_data_1_in_bits),
    .io_data_1_out_valid(PE_48_io_data_1_out_valid),
    .io_data_1_out_bits(PE_48_io_data_1_out_bits),
    .io_data_0_in_valid(PE_48_io_data_0_in_valid),
    .io_data_0_in_bits(PE_48_io_data_0_in_bits),
    .io_data_0_out_valid(PE_48_io_data_0_out_valid),
    .io_data_0_out_bits(PE_48_io_data_0_out_bits)
  );
  PE PE_49 ( // @[pe.scala 184:13]
    .clock(PE_49_clock),
    .reset(PE_49_reset),
    .io_data_2_in_valid(PE_49_io_data_2_in_valid),
    .io_data_2_in_bits(PE_49_io_data_2_in_bits),
    .io_data_2_out_valid(PE_49_io_data_2_out_valid),
    .io_data_2_out_bits(PE_49_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_49_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_49_io_data_2_in_ready),
    .io_data_2_out_ready(PE_49_io_data_2_out_ready),
    .io_data_1_in_valid(PE_49_io_data_1_in_valid),
    .io_data_1_in_bits(PE_49_io_data_1_in_bits),
    .io_data_1_out_valid(PE_49_io_data_1_out_valid),
    .io_data_1_out_bits(PE_49_io_data_1_out_bits),
    .io_data_0_in_valid(PE_49_io_data_0_in_valid),
    .io_data_0_in_bits(PE_49_io_data_0_in_bits),
    .io_data_0_out_valid(PE_49_io_data_0_out_valid),
    .io_data_0_out_bits(PE_49_io_data_0_out_bits)
  );
  PE PE_50 ( // @[pe.scala 184:13]
    .clock(PE_50_clock),
    .reset(PE_50_reset),
    .io_data_2_in_valid(PE_50_io_data_2_in_valid),
    .io_data_2_in_bits(PE_50_io_data_2_in_bits),
    .io_data_2_out_valid(PE_50_io_data_2_out_valid),
    .io_data_2_out_bits(PE_50_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_50_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_50_io_data_2_in_ready),
    .io_data_2_out_ready(PE_50_io_data_2_out_ready),
    .io_data_1_in_valid(PE_50_io_data_1_in_valid),
    .io_data_1_in_bits(PE_50_io_data_1_in_bits),
    .io_data_1_out_valid(PE_50_io_data_1_out_valid),
    .io_data_1_out_bits(PE_50_io_data_1_out_bits),
    .io_data_0_in_valid(PE_50_io_data_0_in_valid),
    .io_data_0_in_bits(PE_50_io_data_0_in_bits),
    .io_data_0_out_valid(PE_50_io_data_0_out_valid),
    .io_data_0_out_bits(PE_50_io_data_0_out_bits)
  );
  PE PE_51 ( // @[pe.scala 184:13]
    .clock(PE_51_clock),
    .reset(PE_51_reset),
    .io_data_2_in_valid(PE_51_io_data_2_in_valid),
    .io_data_2_in_bits(PE_51_io_data_2_in_bits),
    .io_data_2_out_valid(PE_51_io_data_2_out_valid),
    .io_data_2_out_bits(PE_51_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_51_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_51_io_data_2_in_ready),
    .io_data_2_out_ready(PE_51_io_data_2_out_ready),
    .io_data_1_in_valid(PE_51_io_data_1_in_valid),
    .io_data_1_in_bits(PE_51_io_data_1_in_bits),
    .io_data_1_out_valid(PE_51_io_data_1_out_valid),
    .io_data_1_out_bits(PE_51_io_data_1_out_bits),
    .io_data_0_in_valid(PE_51_io_data_0_in_valid),
    .io_data_0_in_bits(PE_51_io_data_0_in_bits),
    .io_data_0_out_valid(PE_51_io_data_0_out_valid),
    .io_data_0_out_bits(PE_51_io_data_0_out_bits)
  );
  PE PE_52 ( // @[pe.scala 184:13]
    .clock(PE_52_clock),
    .reset(PE_52_reset),
    .io_data_2_in_valid(PE_52_io_data_2_in_valid),
    .io_data_2_in_bits(PE_52_io_data_2_in_bits),
    .io_data_2_out_valid(PE_52_io_data_2_out_valid),
    .io_data_2_out_bits(PE_52_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_52_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_52_io_data_2_in_ready),
    .io_data_2_out_ready(PE_52_io_data_2_out_ready),
    .io_data_1_in_valid(PE_52_io_data_1_in_valid),
    .io_data_1_in_bits(PE_52_io_data_1_in_bits),
    .io_data_1_out_valid(PE_52_io_data_1_out_valid),
    .io_data_1_out_bits(PE_52_io_data_1_out_bits),
    .io_data_0_in_valid(PE_52_io_data_0_in_valid),
    .io_data_0_in_bits(PE_52_io_data_0_in_bits),
    .io_data_0_out_valid(PE_52_io_data_0_out_valid),
    .io_data_0_out_bits(PE_52_io_data_0_out_bits)
  );
  PE PE_53 ( // @[pe.scala 184:13]
    .clock(PE_53_clock),
    .reset(PE_53_reset),
    .io_data_2_in_valid(PE_53_io_data_2_in_valid),
    .io_data_2_in_bits(PE_53_io_data_2_in_bits),
    .io_data_2_out_valid(PE_53_io_data_2_out_valid),
    .io_data_2_out_bits(PE_53_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_53_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_53_io_data_2_in_ready),
    .io_data_2_out_ready(PE_53_io_data_2_out_ready),
    .io_data_1_in_valid(PE_53_io_data_1_in_valid),
    .io_data_1_in_bits(PE_53_io_data_1_in_bits),
    .io_data_1_out_valid(PE_53_io_data_1_out_valid),
    .io_data_1_out_bits(PE_53_io_data_1_out_bits),
    .io_data_0_in_valid(PE_53_io_data_0_in_valid),
    .io_data_0_in_bits(PE_53_io_data_0_in_bits),
    .io_data_0_out_valid(PE_53_io_data_0_out_valid),
    .io_data_0_out_bits(PE_53_io_data_0_out_bits)
  );
  PE PE_54 ( // @[pe.scala 184:13]
    .clock(PE_54_clock),
    .reset(PE_54_reset),
    .io_data_2_in_valid(PE_54_io_data_2_in_valid),
    .io_data_2_in_bits(PE_54_io_data_2_in_bits),
    .io_data_2_out_valid(PE_54_io_data_2_out_valid),
    .io_data_2_out_bits(PE_54_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_54_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_54_io_data_2_in_ready),
    .io_data_2_out_ready(PE_54_io_data_2_out_ready),
    .io_data_1_in_valid(PE_54_io_data_1_in_valid),
    .io_data_1_in_bits(PE_54_io_data_1_in_bits),
    .io_data_1_out_valid(PE_54_io_data_1_out_valid),
    .io_data_1_out_bits(PE_54_io_data_1_out_bits),
    .io_data_0_in_valid(PE_54_io_data_0_in_valid),
    .io_data_0_in_bits(PE_54_io_data_0_in_bits),
    .io_data_0_out_valid(PE_54_io_data_0_out_valid),
    .io_data_0_out_bits(PE_54_io_data_0_out_bits)
  );
  PE PE_55 ( // @[pe.scala 184:13]
    .clock(PE_55_clock),
    .reset(PE_55_reset),
    .io_data_2_in_valid(PE_55_io_data_2_in_valid),
    .io_data_2_in_bits(PE_55_io_data_2_in_bits),
    .io_data_2_out_valid(PE_55_io_data_2_out_valid),
    .io_data_2_out_bits(PE_55_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_55_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_55_io_data_2_in_ready),
    .io_data_2_out_ready(PE_55_io_data_2_out_ready),
    .io_data_1_in_valid(PE_55_io_data_1_in_valid),
    .io_data_1_in_bits(PE_55_io_data_1_in_bits),
    .io_data_1_out_valid(PE_55_io_data_1_out_valid),
    .io_data_1_out_bits(PE_55_io_data_1_out_bits),
    .io_data_0_in_valid(PE_55_io_data_0_in_valid),
    .io_data_0_in_bits(PE_55_io_data_0_in_bits),
    .io_data_0_out_valid(PE_55_io_data_0_out_valid),
    .io_data_0_out_bits(PE_55_io_data_0_out_bits)
  );
  PE PE_56 ( // @[pe.scala 184:13]
    .clock(PE_56_clock),
    .reset(PE_56_reset),
    .io_data_2_in_valid(PE_56_io_data_2_in_valid),
    .io_data_2_in_bits(PE_56_io_data_2_in_bits),
    .io_data_2_out_valid(PE_56_io_data_2_out_valid),
    .io_data_2_out_bits(PE_56_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_56_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_56_io_data_2_in_ready),
    .io_data_2_out_ready(PE_56_io_data_2_out_ready),
    .io_data_1_in_valid(PE_56_io_data_1_in_valid),
    .io_data_1_in_bits(PE_56_io_data_1_in_bits),
    .io_data_1_out_valid(PE_56_io_data_1_out_valid),
    .io_data_1_out_bits(PE_56_io_data_1_out_bits),
    .io_data_0_in_valid(PE_56_io_data_0_in_valid),
    .io_data_0_in_bits(PE_56_io_data_0_in_bits),
    .io_data_0_out_valid(PE_56_io_data_0_out_valid),
    .io_data_0_out_bits(PE_56_io_data_0_out_bits)
  );
  PE PE_57 ( // @[pe.scala 184:13]
    .clock(PE_57_clock),
    .reset(PE_57_reset),
    .io_data_2_in_valid(PE_57_io_data_2_in_valid),
    .io_data_2_in_bits(PE_57_io_data_2_in_bits),
    .io_data_2_out_valid(PE_57_io_data_2_out_valid),
    .io_data_2_out_bits(PE_57_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_57_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_57_io_data_2_in_ready),
    .io_data_2_out_ready(PE_57_io_data_2_out_ready),
    .io_data_1_in_valid(PE_57_io_data_1_in_valid),
    .io_data_1_in_bits(PE_57_io_data_1_in_bits),
    .io_data_1_out_valid(PE_57_io_data_1_out_valid),
    .io_data_1_out_bits(PE_57_io_data_1_out_bits),
    .io_data_0_in_valid(PE_57_io_data_0_in_valid),
    .io_data_0_in_bits(PE_57_io_data_0_in_bits),
    .io_data_0_out_valid(PE_57_io_data_0_out_valid),
    .io_data_0_out_bits(PE_57_io_data_0_out_bits)
  );
  PE PE_58 ( // @[pe.scala 184:13]
    .clock(PE_58_clock),
    .reset(PE_58_reset),
    .io_data_2_in_valid(PE_58_io_data_2_in_valid),
    .io_data_2_in_bits(PE_58_io_data_2_in_bits),
    .io_data_2_out_valid(PE_58_io_data_2_out_valid),
    .io_data_2_out_bits(PE_58_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_58_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_58_io_data_2_in_ready),
    .io_data_2_out_ready(PE_58_io_data_2_out_ready),
    .io_data_1_in_valid(PE_58_io_data_1_in_valid),
    .io_data_1_in_bits(PE_58_io_data_1_in_bits),
    .io_data_1_out_valid(PE_58_io_data_1_out_valid),
    .io_data_1_out_bits(PE_58_io_data_1_out_bits),
    .io_data_0_in_valid(PE_58_io_data_0_in_valid),
    .io_data_0_in_bits(PE_58_io_data_0_in_bits),
    .io_data_0_out_valid(PE_58_io_data_0_out_valid),
    .io_data_0_out_bits(PE_58_io_data_0_out_bits)
  );
  PE PE_59 ( // @[pe.scala 184:13]
    .clock(PE_59_clock),
    .reset(PE_59_reset),
    .io_data_2_in_valid(PE_59_io_data_2_in_valid),
    .io_data_2_in_bits(PE_59_io_data_2_in_bits),
    .io_data_2_out_valid(PE_59_io_data_2_out_valid),
    .io_data_2_out_bits(PE_59_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_59_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_59_io_data_2_in_ready),
    .io_data_2_out_ready(PE_59_io_data_2_out_ready),
    .io_data_1_in_valid(PE_59_io_data_1_in_valid),
    .io_data_1_in_bits(PE_59_io_data_1_in_bits),
    .io_data_1_out_valid(PE_59_io_data_1_out_valid),
    .io_data_1_out_bits(PE_59_io_data_1_out_bits),
    .io_data_0_in_valid(PE_59_io_data_0_in_valid),
    .io_data_0_in_bits(PE_59_io_data_0_in_bits),
    .io_data_0_out_valid(PE_59_io_data_0_out_valid),
    .io_data_0_out_bits(PE_59_io_data_0_out_bits)
  );
  PE PE_60 ( // @[pe.scala 184:13]
    .clock(PE_60_clock),
    .reset(PE_60_reset),
    .io_data_2_in_valid(PE_60_io_data_2_in_valid),
    .io_data_2_in_bits(PE_60_io_data_2_in_bits),
    .io_data_2_out_valid(PE_60_io_data_2_out_valid),
    .io_data_2_out_bits(PE_60_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_60_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_60_io_data_2_in_ready),
    .io_data_2_out_ready(PE_60_io_data_2_out_ready),
    .io_data_1_in_valid(PE_60_io_data_1_in_valid),
    .io_data_1_in_bits(PE_60_io_data_1_in_bits),
    .io_data_1_out_valid(PE_60_io_data_1_out_valid),
    .io_data_1_out_bits(PE_60_io_data_1_out_bits),
    .io_data_0_in_valid(PE_60_io_data_0_in_valid),
    .io_data_0_in_bits(PE_60_io_data_0_in_bits),
    .io_data_0_out_valid(PE_60_io_data_0_out_valid),
    .io_data_0_out_bits(PE_60_io_data_0_out_bits)
  );
  PE PE_61 ( // @[pe.scala 184:13]
    .clock(PE_61_clock),
    .reset(PE_61_reset),
    .io_data_2_in_valid(PE_61_io_data_2_in_valid),
    .io_data_2_in_bits(PE_61_io_data_2_in_bits),
    .io_data_2_out_valid(PE_61_io_data_2_out_valid),
    .io_data_2_out_bits(PE_61_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_61_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_61_io_data_2_in_ready),
    .io_data_2_out_ready(PE_61_io_data_2_out_ready),
    .io_data_1_in_valid(PE_61_io_data_1_in_valid),
    .io_data_1_in_bits(PE_61_io_data_1_in_bits),
    .io_data_1_out_valid(PE_61_io_data_1_out_valid),
    .io_data_1_out_bits(PE_61_io_data_1_out_bits),
    .io_data_0_in_valid(PE_61_io_data_0_in_valid),
    .io_data_0_in_bits(PE_61_io_data_0_in_bits),
    .io_data_0_out_valid(PE_61_io_data_0_out_valid),
    .io_data_0_out_bits(PE_61_io_data_0_out_bits)
  );
  PE PE_62 ( // @[pe.scala 184:13]
    .clock(PE_62_clock),
    .reset(PE_62_reset),
    .io_data_2_in_valid(PE_62_io_data_2_in_valid),
    .io_data_2_in_bits(PE_62_io_data_2_in_bits),
    .io_data_2_out_valid(PE_62_io_data_2_out_valid),
    .io_data_2_out_bits(PE_62_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_62_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_62_io_data_2_in_ready),
    .io_data_2_out_ready(PE_62_io_data_2_out_ready),
    .io_data_1_in_valid(PE_62_io_data_1_in_valid),
    .io_data_1_in_bits(PE_62_io_data_1_in_bits),
    .io_data_1_out_valid(PE_62_io_data_1_out_valid),
    .io_data_1_out_bits(PE_62_io_data_1_out_bits),
    .io_data_0_in_valid(PE_62_io_data_0_in_valid),
    .io_data_0_in_bits(PE_62_io_data_0_in_bits),
    .io_data_0_out_valid(PE_62_io_data_0_out_valid),
    .io_data_0_out_bits(PE_62_io_data_0_out_bits)
  );
  PE PE_63 ( // @[pe.scala 184:13]
    .clock(PE_63_clock),
    .reset(PE_63_reset),
    .io_data_2_in_valid(PE_63_io_data_2_in_valid),
    .io_data_2_in_bits(PE_63_io_data_2_in_bits),
    .io_data_2_out_valid(PE_63_io_data_2_out_valid),
    .io_data_2_out_bits(PE_63_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_63_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_63_io_data_2_in_ready),
    .io_data_2_out_ready(PE_63_io_data_2_out_ready),
    .io_data_1_in_valid(PE_63_io_data_1_in_valid),
    .io_data_1_in_bits(PE_63_io_data_1_in_bits),
    .io_data_1_out_valid(PE_63_io_data_1_out_valid),
    .io_data_1_out_bits(PE_63_io_data_1_out_bits),
    .io_data_0_in_valid(PE_63_io_data_0_in_valid),
    .io_data_0_in_bits(PE_63_io_data_0_in_bits),
    .io_data_0_out_valid(PE_63_io_data_0_out_valid),
    .io_data_0_out_bits(PE_63_io_data_0_out_bits)
  );
  PE PE_64 ( // @[pe.scala 184:13]
    .clock(PE_64_clock),
    .reset(PE_64_reset),
    .io_data_2_in_valid(PE_64_io_data_2_in_valid),
    .io_data_2_in_bits(PE_64_io_data_2_in_bits),
    .io_data_2_out_valid(PE_64_io_data_2_out_valid),
    .io_data_2_out_bits(PE_64_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_64_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_64_io_data_2_in_ready),
    .io_data_2_out_ready(PE_64_io_data_2_out_ready),
    .io_data_1_in_valid(PE_64_io_data_1_in_valid),
    .io_data_1_in_bits(PE_64_io_data_1_in_bits),
    .io_data_1_out_valid(PE_64_io_data_1_out_valid),
    .io_data_1_out_bits(PE_64_io_data_1_out_bits),
    .io_data_0_in_valid(PE_64_io_data_0_in_valid),
    .io_data_0_in_bits(PE_64_io_data_0_in_bits),
    .io_data_0_out_valid(PE_64_io_data_0_out_valid),
    .io_data_0_out_bits(PE_64_io_data_0_out_bits)
  );
  PE PE_65 ( // @[pe.scala 184:13]
    .clock(PE_65_clock),
    .reset(PE_65_reset),
    .io_data_2_in_valid(PE_65_io_data_2_in_valid),
    .io_data_2_in_bits(PE_65_io_data_2_in_bits),
    .io_data_2_out_valid(PE_65_io_data_2_out_valid),
    .io_data_2_out_bits(PE_65_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_65_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_65_io_data_2_in_ready),
    .io_data_2_out_ready(PE_65_io_data_2_out_ready),
    .io_data_1_in_valid(PE_65_io_data_1_in_valid),
    .io_data_1_in_bits(PE_65_io_data_1_in_bits),
    .io_data_1_out_valid(PE_65_io_data_1_out_valid),
    .io_data_1_out_bits(PE_65_io_data_1_out_bits),
    .io_data_0_in_valid(PE_65_io_data_0_in_valid),
    .io_data_0_in_bits(PE_65_io_data_0_in_bits),
    .io_data_0_out_valid(PE_65_io_data_0_out_valid),
    .io_data_0_out_bits(PE_65_io_data_0_out_bits)
  );
  PE PE_66 ( // @[pe.scala 184:13]
    .clock(PE_66_clock),
    .reset(PE_66_reset),
    .io_data_2_in_valid(PE_66_io_data_2_in_valid),
    .io_data_2_in_bits(PE_66_io_data_2_in_bits),
    .io_data_2_out_valid(PE_66_io_data_2_out_valid),
    .io_data_2_out_bits(PE_66_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_66_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_66_io_data_2_in_ready),
    .io_data_2_out_ready(PE_66_io_data_2_out_ready),
    .io_data_1_in_valid(PE_66_io_data_1_in_valid),
    .io_data_1_in_bits(PE_66_io_data_1_in_bits),
    .io_data_1_out_valid(PE_66_io_data_1_out_valid),
    .io_data_1_out_bits(PE_66_io_data_1_out_bits),
    .io_data_0_in_valid(PE_66_io_data_0_in_valid),
    .io_data_0_in_bits(PE_66_io_data_0_in_bits),
    .io_data_0_out_valid(PE_66_io_data_0_out_valid),
    .io_data_0_out_bits(PE_66_io_data_0_out_bits)
  );
  PE PE_67 ( // @[pe.scala 184:13]
    .clock(PE_67_clock),
    .reset(PE_67_reset),
    .io_data_2_in_valid(PE_67_io_data_2_in_valid),
    .io_data_2_in_bits(PE_67_io_data_2_in_bits),
    .io_data_2_out_valid(PE_67_io_data_2_out_valid),
    .io_data_2_out_bits(PE_67_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_67_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_67_io_data_2_in_ready),
    .io_data_2_out_ready(PE_67_io_data_2_out_ready),
    .io_data_1_in_valid(PE_67_io_data_1_in_valid),
    .io_data_1_in_bits(PE_67_io_data_1_in_bits),
    .io_data_1_out_valid(PE_67_io_data_1_out_valid),
    .io_data_1_out_bits(PE_67_io_data_1_out_bits),
    .io_data_0_in_valid(PE_67_io_data_0_in_valid),
    .io_data_0_in_bits(PE_67_io_data_0_in_bits),
    .io_data_0_out_valid(PE_67_io_data_0_out_valid),
    .io_data_0_out_bits(PE_67_io_data_0_out_bits)
  );
  PE PE_68 ( // @[pe.scala 184:13]
    .clock(PE_68_clock),
    .reset(PE_68_reset),
    .io_data_2_in_valid(PE_68_io_data_2_in_valid),
    .io_data_2_in_bits(PE_68_io_data_2_in_bits),
    .io_data_2_out_valid(PE_68_io_data_2_out_valid),
    .io_data_2_out_bits(PE_68_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_68_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_68_io_data_2_in_ready),
    .io_data_2_out_ready(PE_68_io_data_2_out_ready),
    .io_data_1_in_valid(PE_68_io_data_1_in_valid),
    .io_data_1_in_bits(PE_68_io_data_1_in_bits),
    .io_data_1_out_valid(PE_68_io_data_1_out_valid),
    .io_data_1_out_bits(PE_68_io_data_1_out_bits),
    .io_data_0_in_valid(PE_68_io_data_0_in_valid),
    .io_data_0_in_bits(PE_68_io_data_0_in_bits),
    .io_data_0_out_valid(PE_68_io_data_0_out_valid),
    .io_data_0_out_bits(PE_68_io_data_0_out_bits)
  );
  PE PE_69 ( // @[pe.scala 184:13]
    .clock(PE_69_clock),
    .reset(PE_69_reset),
    .io_data_2_in_valid(PE_69_io_data_2_in_valid),
    .io_data_2_in_bits(PE_69_io_data_2_in_bits),
    .io_data_2_out_valid(PE_69_io_data_2_out_valid),
    .io_data_2_out_bits(PE_69_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_69_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_69_io_data_2_in_ready),
    .io_data_2_out_ready(PE_69_io_data_2_out_ready),
    .io_data_1_in_valid(PE_69_io_data_1_in_valid),
    .io_data_1_in_bits(PE_69_io_data_1_in_bits),
    .io_data_1_out_valid(PE_69_io_data_1_out_valid),
    .io_data_1_out_bits(PE_69_io_data_1_out_bits),
    .io_data_0_in_valid(PE_69_io_data_0_in_valid),
    .io_data_0_in_bits(PE_69_io_data_0_in_bits),
    .io_data_0_out_valid(PE_69_io_data_0_out_valid),
    .io_data_0_out_bits(PE_69_io_data_0_out_bits)
  );
  PE PE_70 ( // @[pe.scala 184:13]
    .clock(PE_70_clock),
    .reset(PE_70_reset),
    .io_data_2_in_valid(PE_70_io_data_2_in_valid),
    .io_data_2_in_bits(PE_70_io_data_2_in_bits),
    .io_data_2_out_valid(PE_70_io_data_2_out_valid),
    .io_data_2_out_bits(PE_70_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_70_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_70_io_data_2_in_ready),
    .io_data_2_out_ready(PE_70_io_data_2_out_ready),
    .io_data_1_in_valid(PE_70_io_data_1_in_valid),
    .io_data_1_in_bits(PE_70_io_data_1_in_bits),
    .io_data_1_out_valid(PE_70_io_data_1_out_valid),
    .io_data_1_out_bits(PE_70_io_data_1_out_bits),
    .io_data_0_in_valid(PE_70_io_data_0_in_valid),
    .io_data_0_in_bits(PE_70_io_data_0_in_bits),
    .io_data_0_out_valid(PE_70_io_data_0_out_valid),
    .io_data_0_out_bits(PE_70_io_data_0_out_bits)
  );
  PE PE_71 ( // @[pe.scala 184:13]
    .clock(PE_71_clock),
    .reset(PE_71_reset),
    .io_data_2_in_valid(PE_71_io_data_2_in_valid),
    .io_data_2_in_bits(PE_71_io_data_2_in_bits),
    .io_data_2_out_valid(PE_71_io_data_2_out_valid),
    .io_data_2_out_bits(PE_71_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_71_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_71_io_data_2_in_ready),
    .io_data_2_out_ready(PE_71_io_data_2_out_ready),
    .io_data_1_in_valid(PE_71_io_data_1_in_valid),
    .io_data_1_in_bits(PE_71_io_data_1_in_bits),
    .io_data_1_out_valid(PE_71_io_data_1_out_valid),
    .io_data_1_out_bits(PE_71_io_data_1_out_bits),
    .io_data_0_in_valid(PE_71_io_data_0_in_valid),
    .io_data_0_in_bits(PE_71_io_data_0_in_bits),
    .io_data_0_out_valid(PE_71_io_data_0_out_valid),
    .io_data_0_out_bits(PE_71_io_data_0_out_bits)
  );
  PE PE_72 ( // @[pe.scala 184:13]
    .clock(PE_72_clock),
    .reset(PE_72_reset),
    .io_data_2_in_valid(PE_72_io_data_2_in_valid),
    .io_data_2_in_bits(PE_72_io_data_2_in_bits),
    .io_data_2_out_valid(PE_72_io_data_2_out_valid),
    .io_data_2_out_bits(PE_72_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_72_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_72_io_data_2_in_ready),
    .io_data_2_out_ready(PE_72_io_data_2_out_ready),
    .io_data_1_in_valid(PE_72_io_data_1_in_valid),
    .io_data_1_in_bits(PE_72_io_data_1_in_bits),
    .io_data_1_out_valid(PE_72_io_data_1_out_valid),
    .io_data_1_out_bits(PE_72_io_data_1_out_bits),
    .io_data_0_in_valid(PE_72_io_data_0_in_valid),
    .io_data_0_in_bits(PE_72_io_data_0_in_bits),
    .io_data_0_out_valid(PE_72_io_data_0_out_valid),
    .io_data_0_out_bits(PE_72_io_data_0_out_bits)
  );
  PE PE_73 ( // @[pe.scala 184:13]
    .clock(PE_73_clock),
    .reset(PE_73_reset),
    .io_data_2_in_valid(PE_73_io_data_2_in_valid),
    .io_data_2_in_bits(PE_73_io_data_2_in_bits),
    .io_data_2_out_valid(PE_73_io_data_2_out_valid),
    .io_data_2_out_bits(PE_73_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_73_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_73_io_data_2_in_ready),
    .io_data_2_out_ready(PE_73_io_data_2_out_ready),
    .io_data_1_in_valid(PE_73_io_data_1_in_valid),
    .io_data_1_in_bits(PE_73_io_data_1_in_bits),
    .io_data_1_out_valid(PE_73_io_data_1_out_valid),
    .io_data_1_out_bits(PE_73_io_data_1_out_bits),
    .io_data_0_in_valid(PE_73_io_data_0_in_valid),
    .io_data_0_in_bits(PE_73_io_data_0_in_bits),
    .io_data_0_out_valid(PE_73_io_data_0_out_valid),
    .io_data_0_out_bits(PE_73_io_data_0_out_bits)
  );
  PE PE_74 ( // @[pe.scala 184:13]
    .clock(PE_74_clock),
    .reset(PE_74_reset),
    .io_data_2_in_valid(PE_74_io_data_2_in_valid),
    .io_data_2_in_bits(PE_74_io_data_2_in_bits),
    .io_data_2_out_valid(PE_74_io_data_2_out_valid),
    .io_data_2_out_bits(PE_74_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_74_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_74_io_data_2_in_ready),
    .io_data_2_out_ready(PE_74_io_data_2_out_ready),
    .io_data_1_in_valid(PE_74_io_data_1_in_valid),
    .io_data_1_in_bits(PE_74_io_data_1_in_bits),
    .io_data_1_out_valid(PE_74_io_data_1_out_valid),
    .io_data_1_out_bits(PE_74_io_data_1_out_bits),
    .io_data_0_in_valid(PE_74_io_data_0_in_valid),
    .io_data_0_in_bits(PE_74_io_data_0_in_bits),
    .io_data_0_out_valid(PE_74_io_data_0_out_valid),
    .io_data_0_out_bits(PE_74_io_data_0_out_bits)
  );
  PE PE_75 ( // @[pe.scala 184:13]
    .clock(PE_75_clock),
    .reset(PE_75_reset),
    .io_data_2_in_valid(PE_75_io_data_2_in_valid),
    .io_data_2_in_bits(PE_75_io_data_2_in_bits),
    .io_data_2_out_valid(PE_75_io_data_2_out_valid),
    .io_data_2_out_bits(PE_75_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_75_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_75_io_data_2_in_ready),
    .io_data_2_out_ready(PE_75_io_data_2_out_ready),
    .io_data_1_in_valid(PE_75_io_data_1_in_valid),
    .io_data_1_in_bits(PE_75_io_data_1_in_bits),
    .io_data_1_out_valid(PE_75_io_data_1_out_valid),
    .io_data_1_out_bits(PE_75_io_data_1_out_bits),
    .io_data_0_in_valid(PE_75_io_data_0_in_valid),
    .io_data_0_in_bits(PE_75_io_data_0_in_bits),
    .io_data_0_out_valid(PE_75_io_data_0_out_valid),
    .io_data_0_out_bits(PE_75_io_data_0_out_bits)
  );
  PE PE_76 ( // @[pe.scala 184:13]
    .clock(PE_76_clock),
    .reset(PE_76_reset),
    .io_data_2_in_valid(PE_76_io_data_2_in_valid),
    .io_data_2_in_bits(PE_76_io_data_2_in_bits),
    .io_data_2_out_valid(PE_76_io_data_2_out_valid),
    .io_data_2_out_bits(PE_76_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_76_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_76_io_data_2_in_ready),
    .io_data_2_out_ready(PE_76_io_data_2_out_ready),
    .io_data_1_in_valid(PE_76_io_data_1_in_valid),
    .io_data_1_in_bits(PE_76_io_data_1_in_bits),
    .io_data_1_out_valid(PE_76_io_data_1_out_valid),
    .io_data_1_out_bits(PE_76_io_data_1_out_bits),
    .io_data_0_in_valid(PE_76_io_data_0_in_valid),
    .io_data_0_in_bits(PE_76_io_data_0_in_bits),
    .io_data_0_out_valid(PE_76_io_data_0_out_valid),
    .io_data_0_out_bits(PE_76_io_data_0_out_bits)
  );
  PE PE_77 ( // @[pe.scala 184:13]
    .clock(PE_77_clock),
    .reset(PE_77_reset),
    .io_data_2_in_valid(PE_77_io_data_2_in_valid),
    .io_data_2_in_bits(PE_77_io_data_2_in_bits),
    .io_data_2_out_valid(PE_77_io_data_2_out_valid),
    .io_data_2_out_bits(PE_77_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_77_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_77_io_data_2_in_ready),
    .io_data_2_out_ready(PE_77_io_data_2_out_ready),
    .io_data_1_in_valid(PE_77_io_data_1_in_valid),
    .io_data_1_in_bits(PE_77_io_data_1_in_bits),
    .io_data_1_out_valid(PE_77_io_data_1_out_valid),
    .io_data_1_out_bits(PE_77_io_data_1_out_bits),
    .io_data_0_in_valid(PE_77_io_data_0_in_valid),
    .io_data_0_in_bits(PE_77_io_data_0_in_bits),
    .io_data_0_out_valid(PE_77_io_data_0_out_valid),
    .io_data_0_out_bits(PE_77_io_data_0_out_bits)
  );
  PE PE_78 ( // @[pe.scala 184:13]
    .clock(PE_78_clock),
    .reset(PE_78_reset),
    .io_data_2_in_valid(PE_78_io_data_2_in_valid),
    .io_data_2_in_bits(PE_78_io_data_2_in_bits),
    .io_data_2_out_valid(PE_78_io_data_2_out_valid),
    .io_data_2_out_bits(PE_78_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_78_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_78_io_data_2_in_ready),
    .io_data_2_out_ready(PE_78_io_data_2_out_ready),
    .io_data_1_in_valid(PE_78_io_data_1_in_valid),
    .io_data_1_in_bits(PE_78_io_data_1_in_bits),
    .io_data_1_out_valid(PE_78_io_data_1_out_valid),
    .io_data_1_out_bits(PE_78_io_data_1_out_bits),
    .io_data_0_in_valid(PE_78_io_data_0_in_valid),
    .io_data_0_in_bits(PE_78_io_data_0_in_bits),
    .io_data_0_out_valid(PE_78_io_data_0_out_valid),
    .io_data_0_out_bits(PE_78_io_data_0_out_bits)
  );
  PE PE_79 ( // @[pe.scala 184:13]
    .clock(PE_79_clock),
    .reset(PE_79_reset),
    .io_data_2_in_valid(PE_79_io_data_2_in_valid),
    .io_data_2_in_bits(PE_79_io_data_2_in_bits),
    .io_data_2_out_valid(PE_79_io_data_2_out_valid),
    .io_data_2_out_bits(PE_79_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_79_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_79_io_data_2_in_ready),
    .io_data_2_out_ready(PE_79_io_data_2_out_ready),
    .io_data_1_in_valid(PE_79_io_data_1_in_valid),
    .io_data_1_in_bits(PE_79_io_data_1_in_bits),
    .io_data_1_out_valid(PE_79_io_data_1_out_valid),
    .io_data_1_out_bits(PE_79_io_data_1_out_bits),
    .io_data_0_in_valid(PE_79_io_data_0_in_valid),
    .io_data_0_in_bits(PE_79_io_data_0_in_bits),
    .io_data_0_out_valid(PE_79_io_data_0_out_valid),
    .io_data_0_out_bits(PE_79_io_data_0_out_bits)
  );
  PE PE_80 ( // @[pe.scala 184:13]
    .clock(PE_80_clock),
    .reset(PE_80_reset),
    .io_data_2_in_valid(PE_80_io_data_2_in_valid),
    .io_data_2_in_bits(PE_80_io_data_2_in_bits),
    .io_data_2_out_valid(PE_80_io_data_2_out_valid),
    .io_data_2_out_bits(PE_80_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_80_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_80_io_data_2_in_ready),
    .io_data_2_out_ready(PE_80_io_data_2_out_ready),
    .io_data_1_in_valid(PE_80_io_data_1_in_valid),
    .io_data_1_in_bits(PE_80_io_data_1_in_bits),
    .io_data_1_out_valid(PE_80_io_data_1_out_valid),
    .io_data_1_out_bits(PE_80_io_data_1_out_bits),
    .io_data_0_in_valid(PE_80_io_data_0_in_valid),
    .io_data_0_in_bits(PE_80_io_data_0_in_bits),
    .io_data_0_out_valid(PE_80_io_data_0_out_valid),
    .io_data_0_out_bits(PE_80_io_data_0_out_bits)
  );
  PE PE_81 ( // @[pe.scala 184:13]
    .clock(PE_81_clock),
    .reset(PE_81_reset),
    .io_data_2_in_valid(PE_81_io_data_2_in_valid),
    .io_data_2_in_bits(PE_81_io_data_2_in_bits),
    .io_data_2_out_valid(PE_81_io_data_2_out_valid),
    .io_data_2_out_bits(PE_81_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_81_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_81_io_data_2_in_ready),
    .io_data_2_out_ready(PE_81_io_data_2_out_ready),
    .io_data_1_in_valid(PE_81_io_data_1_in_valid),
    .io_data_1_in_bits(PE_81_io_data_1_in_bits),
    .io_data_1_out_valid(PE_81_io_data_1_out_valid),
    .io_data_1_out_bits(PE_81_io_data_1_out_bits),
    .io_data_0_in_valid(PE_81_io_data_0_in_valid),
    .io_data_0_in_bits(PE_81_io_data_0_in_bits),
    .io_data_0_out_valid(PE_81_io_data_0_out_valid),
    .io_data_0_out_bits(PE_81_io_data_0_out_bits)
  );
  PE PE_82 ( // @[pe.scala 184:13]
    .clock(PE_82_clock),
    .reset(PE_82_reset),
    .io_data_2_in_valid(PE_82_io_data_2_in_valid),
    .io_data_2_in_bits(PE_82_io_data_2_in_bits),
    .io_data_2_out_valid(PE_82_io_data_2_out_valid),
    .io_data_2_out_bits(PE_82_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_82_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_82_io_data_2_in_ready),
    .io_data_2_out_ready(PE_82_io_data_2_out_ready),
    .io_data_1_in_valid(PE_82_io_data_1_in_valid),
    .io_data_1_in_bits(PE_82_io_data_1_in_bits),
    .io_data_1_out_valid(PE_82_io_data_1_out_valid),
    .io_data_1_out_bits(PE_82_io_data_1_out_bits),
    .io_data_0_in_valid(PE_82_io_data_0_in_valid),
    .io_data_0_in_bits(PE_82_io_data_0_in_bits),
    .io_data_0_out_valid(PE_82_io_data_0_out_valid),
    .io_data_0_out_bits(PE_82_io_data_0_out_bits)
  );
  PE PE_83 ( // @[pe.scala 184:13]
    .clock(PE_83_clock),
    .reset(PE_83_reset),
    .io_data_2_in_valid(PE_83_io_data_2_in_valid),
    .io_data_2_in_bits(PE_83_io_data_2_in_bits),
    .io_data_2_out_valid(PE_83_io_data_2_out_valid),
    .io_data_2_out_bits(PE_83_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_83_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_83_io_data_2_in_ready),
    .io_data_2_out_ready(PE_83_io_data_2_out_ready),
    .io_data_1_in_valid(PE_83_io_data_1_in_valid),
    .io_data_1_in_bits(PE_83_io_data_1_in_bits),
    .io_data_1_out_valid(PE_83_io_data_1_out_valid),
    .io_data_1_out_bits(PE_83_io_data_1_out_bits),
    .io_data_0_in_valid(PE_83_io_data_0_in_valid),
    .io_data_0_in_bits(PE_83_io_data_0_in_bits),
    .io_data_0_out_valid(PE_83_io_data_0_out_valid),
    .io_data_0_out_bits(PE_83_io_data_0_out_bits)
  );
  PE PE_84 ( // @[pe.scala 184:13]
    .clock(PE_84_clock),
    .reset(PE_84_reset),
    .io_data_2_in_valid(PE_84_io_data_2_in_valid),
    .io_data_2_in_bits(PE_84_io_data_2_in_bits),
    .io_data_2_out_valid(PE_84_io_data_2_out_valid),
    .io_data_2_out_bits(PE_84_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_84_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_84_io_data_2_in_ready),
    .io_data_2_out_ready(PE_84_io_data_2_out_ready),
    .io_data_1_in_valid(PE_84_io_data_1_in_valid),
    .io_data_1_in_bits(PE_84_io_data_1_in_bits),
    .io_data_1_out_valid(PE_84_io_data_1_out_valid),
    .io_data_1_out_bits(PE_84_io_data_1_out_bits),
    .io_data_0_in_valid(PE_84_io_data_0_in_valid),
    .io_data_0_in_bits(PE_84_io_data_0_in_bits),
    .io_data_0_out_valid(PE_84_io_data_0_out_valid),
    .io_data_0_out_bits(PE_84_io_data_0_out_bits)
  );
  PE PE_85 ( // @[pe.scala 184:13]
    .clock(PE_85_clock),
    .reset(PE_85_reset),
    .io_data_2_in_valid(PE_85_io_data_2_in_valid),
    .io_data_2_in_bits(PE_85_io_data_2_in_bits),
    .io_data_2_out_valid(PE_85_io_data_2_out_valid),
    .io_data_2_out_bits(PE_85_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_85_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_85_io_data_2_in_ready),
    .io_data_2_out_ready(PE_85_io_data_2_out_ready),
    .io_data_1_in_valid(PE_85_io_data_1_in_valid),
    .io_data_1_in_bits(PE_85_io_data_1_in_bits),
    .io_data_1_out_valid(PE_85_io_data_1_out_valid),
    .io_data_1_out_bits(PE_85_io_data_1_out_bits),
    .io_data_0_in_valid(PE_85_io_data_0_in_valid),
    .io_data_0_in_bits(PE_85_io_data_0_in_bits),
    .io_data_0_out_valid(PE_85_io_data_0_out_valid),
    .io_data_0_out_bits(PE_85_io_data_0_out_bits)
  );
  PE PE_86 ( // @[pe.scala 184:13]
    .clock(PE_86_clock),
    .reset(PE_86_reset),
    .io_data_2_in_valid(PE_86_io_data_2_in_valid),
    .io_data_2_in_bits(PE_86_io_data_2_in_bits),
    .io_data_2_out_valid(PE_86_io_data_2_out_valid),
    .io_data_2_out_bits(PE_86_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_86_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_86_io_data_2_in_ready),
    .io_data_2_out_ready(PE_86_io_data_2_out_ready),
    .io_data_1_in_valid(PE_86_io_data_1_in_valid),
    .io_data_1_in_bits(PE_86_io_data_1_in_bits),
    .io_data_1_out_valid(PE_86_io_data_1_out_valid),
    .io_data_1_out_bits(PE_86_io_data_1_out_bits),
    .io_data_0_in_valid(PE_86_io_data_0_in_valid),
    .io_data_0_in_bits(PE_86_io_data_0_in_bits),
    .io_data_0_out_valid(PE_86_io_data_0_out_valid),
    .io_data_0_out_bits(PE_86_io_data_0_out_bits)
  );
  PE PE_87 ( // @[pe.scala 184:13]
    .clock(PE_87_clock),
    .reset(PE_87_reset),
    .io_data_2_in_valid(PE_87_io_data_2_in_valid),
    .io_data_2_in_bits(PE_87_io_data_2_in_bits),
    .io_data_2_out_valid(PE_87_io_data_2_out_valid),
    .io_data_2_out_bits(PE_87_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_87_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_87_io_data_2_in_ready),
    .io_data_2_out_ready(PE_87_io_data_2_out_ready),
    .io_data_1_in_valid(PE_87_io_data_1_in_valid),
    .io_data_1_in_bits(PE_87_io_data_1_in_bits),
    .io_data_1_out_valid(PE_87_io_data_1_out_valid),
    .io_data_1_out_bits(PE_87_io_data_1_out_bits),
    .io_data_0_in_valid(PE_87_io_data_0_in_valid),
    .io_data_0_in_bits(PE_87_io_data_0_in_bits),
    .io_data_0_out_valid(PE_87_io_data_0_out_valid),
    .io_data_0_out_bits(PE_87_io_data_0_out_bits)
  );
  PE PE_88 ( // @[pe.scala 184:13]
    .clock(PE_88_clock),
    .reset(PE_88_reset),
    .io_data_2_in_valid(PE_88_io_data_2_in_valid),
    .io_data_2_in_bits(PE_88_io_data_2_in_bits),
    .io_data_2_out_valid(PE_88_io_data_2_out_valid),
    .io_data_2_out_bits(PE_88_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_88_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_88_io_data_2_in_ready),
    .io_data_2_out_ready(PE_88_io_data_2_out_ready),
    .io_data_1_in_valid(PE_88_io_data_1_in_valid),
    .io_data_1_in_bits(PE_88_io_data_1_in_bits),
    .io_data_1_out_valid(PE_88_io_data_1_out_valid),
    .io_data_1_out_bits(PE_88_io_data_1_out_bits),
    .io_data_0_in_valid(PE_88_io_data_0_in_valid),
    .io_data_0_in_bits(PE_88_io_data_0_in_bits),
    .io_data_0_out_valid(PE_88_io_data_0_out_valid),
    .io_data_0_out_bits(PE_88_io_data_0_out_bits)
  );
  PE PE_89 ( // @[pe.scala 184:13]
    .clock(PE_89_clock),
    .reset(PE_89_reset),
    .io_data_2_in_valid(PE_89_io_data_2_in_valid),
    .io_data_2_in_bits(PE_89_io_data_2_in_bits),
    .io_data_2_out_valid(PE_89_io_data_2_out_valid),
    .io_data_2_out_bits(PE_89_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_89_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_89_io_data_2_in_ready),
    .io_data_2_out_ready(PE_89_io_data_2_out_ready),
    .io_data_1_in_valid(PE_89_io_data_1_in_valid),
    .io_data_1_in_bits(PE_89_io_data_1_in_bits),
    .io_data_1_out_valid(PE_89_io_data_1_out_valid),
    .io_data_1_out_bits(PE_89_io_data_1_out_bits),
    .io_data_0_in_valid(PE_89_io_data_0_in_valid),
    .io_data_0_in_bits(PE_89_io_data_0_in_bits),
    .io_data_0_out_valid(PE_89_io_data_0_out_valid),
    .io_data_0_out_bits(PE_89_io_data_0_out_bits)
  );
  PE PE_90 ( // @[pe.scala 184:13]
    .clock(PE_90_clock),
    .reset(PE_90_reset),
    .io_data_2_in_valid(PE_90_io_data_2_in_valid),
    .io_data_2_in_bits(PE_90_io_data_2_in_bits),
    .io_data_2_out_valid(PE_90_io_data_2_out_valid),
    .io_data_2_out_bits(PE_90_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_90_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_90_io_data_2_in_ready),
    .io_data_2_out_ready(PE_90_io_data_2_out_ready),
    .io_data_1_in_valid(PE_90_io_data_1_in_valid),
    .io_data_1_in_bits(PE_90_io_data_1_in_bits),
    .io_data_1_out_valid(PE_90_io_data_1_out_valid),
    .io_data_1_out_bits(PE_90_io_data_1_out_bits),
    .io_data_0_in_valid(PE_90_io_data_0_in_valid),
    .io_data_0_in_bits(PE_90_io_data_0_in_bits),
    .io_data_0_out_valid(PE_90_io_data_0_out_valid),
    .io_data_0_out_bits(PE_90_io_data_0_out_bits)
  );
  PE PE_91 ( // @[pe.scala 184:13]
    .clock(PE_91_clock),
    .reset(PE_91_reset),
    .io_data_2_in_valid(PE_91_io_data_2_in_valid),
    .io_data_2_in_bits(PE_91_io_data_2_in_bits),
    .io_data_2_out_valid(PE_91_io_data_2_out_valid),
    .io_data_2_out_bits(PE_91_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_91_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_91_io_data_2_in_ready),
    .io_data_2_out_ready(PE_91_io_data_2_out_ready),
    .io_data_1_in_valid(PE_91_io_data_1_in_valid),
    .io_data_1_in_bits(PE_91_io_data_1_in_bits),
    .io_data_1_out_valid(PE_91_io_data_1_out_valid),
    .io_data_1_out_bits(PE_91_io_data_1_out_bits),
    .io_data_0_in_valid(PE_91_io_data_0_in_valid),
    .io_data_0_in_bits(PE_91_io_data_0_in_bits),
    .io_data_0_out_valid(PE_91_io_data_0_out_valid),
    .io_data_0_out_bits(PE_91_io_data_0_out_bits)
  );
  PE PE_92 ( // @[pe.scala 184:13]
    .clock(PE_92_clock),
    .reset(PE_92_reset),
    .io_data_2_in_valid(PE_92_io_data_2_in_valid),
    .io_data_2_in_bits(PE_92_io_data_2_in_bits),
    .io_data_2_out_valid(PE_92_io_data_2_out_valid),
    .io_data_2_out_bits(PE_92_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_92_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_92_io_data_2_in_ready),
    .io_data_2_out_ready(PE_92_io_data_2_out_ready),
    .io_data_1_in_valid(PE_92_io_data_1_in_valid),
    .io_data_1_in_bits(PE_92_io_data_1_in_bits),
    .io_data_1_out_valid(PE_92_io_data_1_out_valid),
    .io_data_1_out_bits(PE_92_io_data_1_out_bits),
    .io_data_0_in_valid(PE_92_io_data_0_in_valid),
    .io_data_0_in_bits(PE_92_io_data_0_in_bits),
    .io_data_0_out_valid(PE_92_io_data_0_out_valid),
    .io_data_0_out_bits(PE_92_io_data_0_out_bits)
  );
  PE PE_93 ( // @[pe.scala 184:13]
    .clock(PE_93_clock),
    .reset(PE_93_reset),
    .io_data_2_in_valid(PE_93_io_data_2_in_valid),
    .io_data_2_in_bits(PE_93_io_data_2_in_bits),
    .io_data_2_out_valid(PE_93_io_data_2_out_valid),
    .io_data_2_out_bits(PE_93_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_93_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_93_io_data_2_in_ready),
    .io_data_2_out_ready(PE_93_io_data_2_out_ready),
    .io_data_1_in_valid(PE_93_io_data_1_in_valid),
    .io_data_1_in_bits(PE_93_io_data_1_in_bits),
    .io_data_1_out_valid(PE_93_io_data_1_out_valid),
    .io_data_1_out_bits(PE_93_io_data_1_out_bits),
    .io_data_0_in_valid(PE_93_io_data_0_in_valid),
    .io_data_0_in_bits(PE_93_io_data_0_in_bits),
    .io_data_0_out_valid(PE_93_io_data_0_out_valid),
    .io_data_0_out_bits(PE_93_io_data_0_out_bits)
  );
  PE PE_94 ( // @[pe.scala 184:13]
    .clock(PE_94_clock),
    .reset(PE_94_reset),
    .io_data_2_in_valid(PE_94_io_data_2_in_valid),
    .io_data_2_in_bits(PE_94_io_data_2_in_bits),
    .io_data_2_out_valid(PE_94_io_data_2_out_valid),
    .io_data_2_out_bits(PE_94_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_94_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_94_io_data_2_in_ready),
    .io_data_2_out_ready(PE_94_io_data_2_out_ready),
    .io_data_1_in_valid(PE_94_io_data_1_in_valid),
    .io_data_1_in_bits(PE_94_io_data_1_in_bits),
    .io_data_1_out_valid(PE_94_io_data_1_out_valid),
    .io_data_1_out_bits(PE_94_io_data_1_out_bits),
    .io_data_0_in_valid(PE_94_io_data_0_in_valid),
    .io_data_0_in_bits(PE_94_io_data_0_in_bits),
    .io_data_0_out_valid(PE_94_io_data_0_out_valid),
    .io_data_0_out_bits(PE_94_io_data_0_out_bits)
  );
  PE PE_95 ( // @[pe.scala 184:13]
    .clock(PE_95_clock),
    .reset(PE_95_reset),
    .io_data_2_in_valid(PE_95_io_data_2_in_valid),
    .io_data_2_in_bits(PE_95_io_data_2_in_bits),
    .io_data_2_out_valid(PE_95_io_data_2_out_valid),
    .io_data_2_out_bits(PE_95_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_95_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_95_io_data_2_in_ready),
    .io_data_2_out_ready(PE_95_io_data_2_out_ready),
    .io_data_1_in_valid(PE_95_io_data_1_in_valid),
    .io_data_1_in_bits(PE_95_io_data_1_in_bits),
    .io_data_1_out_valid(PE_95_io_data_1_out_valid),
    .io_data_1_out_bits(PE_95_io_data_1_out_bits),
    .io_data_0_in_valid(PE_95_io_data_0_in_valid),
    .io_data_0_in_bits(PE_95_io_data_0_in_bits),
    .io_data_0_out_valid(PE_95_io_data_0_out_valid),
    .io_data_0_out_bits(PE_95_io_data_0_out_bits)
  );
  PE PE_96 ( // @[pe.scala 184:13]
    .clock(PE_96_clock),
    .reset(PE_96_reset),
    .io_data_2_in_valid(PE_96_io_data_2_in_valid),
    .io_data_2_in_bits(PE_96_io_data_2_in_bits),
    .io_data_2_out_valid(PE_96_io_data_2_out_valid),
    .io_data_2_out_bits(PE_96_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_96_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_96_io_data_2_in_ready),
    .io_data_2_out_ready(PE_96_io_data_2_out_ready),
    .io_data_1_in_valid(PE_96_io_data_1_in_valid),
    .io_data_1_in_bits(PE_96_io_data_1_in_bits),
    .io_data_1_out_valid(PE_96_io_data_1_out_valid),
    .io_data_1_out_bits(PE_96_io_data_1_out_bits),
    .io_data_0_in_valid(PE_96_io_data_0_in_valid),
    .io_data_0_in_bits(PE_96_io_data_0_in_bits),
    .io_data_0_out_valid(PE_96_io_data_0_out_valid),
    .io_data_0_out_bits(PE_96_io_data_0_out_bits)
  );
  PE PE_97 ( // @[pe.scala 184:13]
    .clock(PE_97_clock),
    .reset(PE_97_reset),
    .io_data_2_in_valid(PE_97_io_data_2_in_valid),
    .io_data_2_in_bits(PE_97_io_data_2_in_bits),
    .io_data_2_out_valid(PE_97_io_data_2_out_valid),
    .io_data_2_out_bits(PE_97_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_97_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_97_io_data_2_in_ready),
    .io_data_2_out_ready(PE_97_io_data_2_out_ready),
    .io_data_1_in_valid(PE_97_io_data_1_in_valid),
    .io_data_1_in_bits(PE_97_io_data_1_in_bits),
    .io_data_1_out_valid(PE_97_io_data_1_out_valid),
    .io_data_1_out_bits(PE_97_io_data_1_out_bits),
    .io_data_0_in_valid(PE_97_io_data_0_in_valid),
    .io_data_0_in_bits(PE_97_io_data_0_in_bits),
    .io_data_0_out_valid(PE_97_io_data_0_out_valid),
    .io_data_0_out_bits(PE_97_io_data_0_out_bits)
  );
  PE PE_98 ( // @[pe.scala 184:13]
    .clock(PE_98_clock),
    .reset(PE_98_reset),
    .io_data_2_in_valid(PE_98_io_data_2_in_valid),
    .io_data_2_in_bits(PE_98_io_data_2_in_bits),
    .io_data_2_out_valid(PE_98_io_data_2_out_valid),
    .io_data_2_out_bits(PE_98_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_98_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_98_io_data_2_in_ready),
    .io_data_2_out_ready(PE_98_io_data_2_out_ready),
    .io_data_1_in_valid(PE_98_io_data_1_in_valid),
    .io_data_1_in_bits(PE_98_io_data_1_in_bits),
    .io_data_1_out_valid(PE_98_io_data_1_out_valid),
    .io_data_1_out_bits(PE_98_io_data_1_out_bits),
    .io_data_0_in_valid(PE_98_io_data_0_in_valid),
    .io_data_0_in_bits(PE_98_io_data_0_in_bits),
    .io_data_0_out_valid(PE_98_io_data_0_out_valid),
    .io_data_0_out_bits(PE_98_io_data_0_out_bits)
  );
  PE PE_99 ( // @[pe.scala 184:13]
    .clock(PE_99_clock),
    .reset(PE_99_reset),
    .io_data_2_in_valid(PE_99_io_data_2_in_valid),
    .io_data_2_in_bits(PE_99_io_data_2_in_bits),
    .io_data_2_out_valid(PE_99_io_data_2_out_valid),
    .io_data_2_out_bits(PE_99_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_99_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_99_io_data_2_in_ready),
    .io_data_2_out_ready(PE_99_io_data_2_out_ready),
    .io_data_1_in_valid(PE_99_io_data_1_in_valid),
    .io_data_1_in_bits(PE_99_io_data_1_in_bits),
    .io_data_1_out_valid(PE_99_io_data_1_out_valid),
    .io_data_1_out_bits(PE_99_io_data_1_out_bits),
    .io_data_0_in_valid(PE_99_io_data_0_in_valid),
    .io_data_0_in_bits(PE_99_io_data_0_in_bits),
    .io_data_0_out_valid(PE_99_io_data_0_out_valid),
    .io_data_0_out_bits(PE_99_io_data_0_out_bits)
  );
  PE PE_100 ( // @[pe.scala 184:13]
    .clock(PE_100_clock),
    .reset(PE_100_reset),
    .io_data_2_in_valid(PE_100_io_data_2_in_valid),
    .io_data_2_in_bits(PE_100_io_data_2_in_bits),
    .io_data_2_out_valid(PE_100_io_data_2_out_valid),
    .io_data_2_out_bits(PE_100_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_100_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_100_io_data_2_in_ready),
    .io_data_2_out_ready(PE_100_io_data_2_out_ready),
    .io_data_1_in_valid(PE_100_io_data_1_in_valid),
    .io_data_1_in_bits(PE_100_io_data_1_in_bits),
    .io_data_1_out_valid(PE_100_io_data_1_out_valid),
    .io_data_1_out_bits(PE_100_io_data_1_out_bits),
    .io_data_0_in_valid(PE_100_io_data_0_in_valid),
    .io_data_0_in_bits(PE_100_io_data_0_in_bits),
    .io_data_0_out_valid(PE_100_io_data_0_out_valid),
    .io_data_0_out_bits(PE_100_io_data_0_out_bits)
  );
  PE PE_101 ( // @[pe.scala 184:13]
    .clock(PE_101_clock),
    .reset(PE_101_reset),
    .io_data_2_in_valid(PE_101_io_data_2_in_valid),
    .io_data_2_in_bits(PE_101_io_data_2_in_bits),
    .io_data_2_out_valid(PE_101_io_data_2_out_valid),
    .io_data_2_out_bits(PE_101_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_101_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_101_io_data_2_in_ready),
    .io_data_2_out_ready(PE_101_io_data_2_out_ready),
    .io_data_1_in_valid(PE_101_io_data_1_in_valid),
    .io_data_1_in_bits(PE_101_io_data_1_in_bits),
    .io_data_1_out_valid(PE_101_io_data_1_out_valid),
    .io_data_1_out_bits(PE_101_io_data_1_out_bits),
    .io_data_0_in_valid(PE_101_io_data_0_in_valid),
    .io_data_0_in_bits(PE_101_io_data_0_in_bits),
    .io_data_0_out_valid(PE_101_io_data_0_out_valid),
    .io_data_0_out_bits(PE_101_io_data_0_out_bits)
  );
  PE PE_102 ( // @[pe.scala 184:13]
    .clock(PE_102_clock),
    .reset(PE_102_reset),
    .io_data_2_in_valid(PE_102_io_data_2_in_valid),
    .io_data_2_in_bits(PE_102_io_data_2_in_bits),
    .io_data_2_out_valid(PE_102_io_data_2_out_valid),
    .io_data_2_out_bits(PE_102_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_102_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_102_io_data_2_in_ready),
    .io_data_2_out_ready(PE_102_io_data_2_out_ready),
    .io_data_1_in_valid(PE_102_io_data_1_in_valid),
    .io_data_1_in_bits(PE_102_io_data_1_in_bits),
    .io_data_1_out_valid(PE_102_io_data_1_out_valid),
    .io_data_1_out_bits(PE_102_io_data_1_out_bits),
    .io_data_0_in_valid(PE_102_io_data_0_in_valid),
    .io_data_0_in_bits(PE_102_io_data_0_in_bits),
    .io_data_0_out_valid(PE_102_io_data_0_out_valid),
    .io_data_0_out_bits(PE_102_io_data_0_out_bits)
  );
  PE PE_103 ( // @[pe.scala 184:13]
    .clock(PE_103_clock),
    .reset(PE_103_reset),
    .io_data_2_in_valid(PE_103_io_data_2_in_valid),
    .io_data_2_in_bits(PE_103_io_data_2_in_bits),
    .io_data_2_out_valid(PE_103_io_data_2_out_valid),
    .io_data_2_out_bits(PE_103_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_103_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_103_io_data_2_in_ready),
    .io_data_2_out_ready(PE_103_io_data_2_out_ready),
    .io_data_1_in_valid(PE_103_io_data_1_in_valid),
    .io_data_1_in_bits(PE_103_io_data_1_in_bits),
    .io_data_1_out_valid(PE_103_io_data_1_out_valid),
    .io_data_1_out_bits(PE_103_io_data_1_out_bits),
    .io_data_0_in_valid(PE_103_io_data_0_in_valid),
    .io_data_0_in_bits(PE_103_io_data_0_in_bits),
    .io_data_0_out_valid(PE_103_io_data_0_out_valid),
    .io_data_0_out_bits(PE_103_io_data_0_out_bits)
  );
  PE PE_104 ( // @[pe.scala 184:13]
    .clock(PE_104_clock),
    .reset(PE_104_reset),
    .io_data_2_in_valid(PE_104_io_data_2_in_valid),
    .io_data_2_in_bits(PE_104_io_data_2_in_bits),
    .io_data_2_out_valid(PE_104_io_data_2_out_valid),
    .io_data_2_out_bits(PE_104_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_104_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_104_io_data_2_in_ready),
    .io_data_2_out_ready(PE_104_io_data_2_out_ready),
    .io_data_1_in_valid(PE_104_io_data_1_in_valid),
    .io_data_1_in_bits(PE_104_io_data_1_in_bits),
    .io_data_1_out_valid(PE_104_io_data_1_out_valid),
    .io_data_1_out_bits(PE_104_io_data_1_out_bits),
    .io_data_0_in_valid(PE_104_io_data_0_in_valid),
    .io_data_0_in_bits(PE_104_io_data_0_in_bits),
    .io_data_0_out_valid(PE_104_io_data_0_out_valid),
    .io_data_0_out_bits(PE_104_io_data_0_out_bits)
  );
  PE PE_105 ( // @[pe.scala 184:13]
    .clock(PE_105_clock),
    .reset(PE_105_reset),
    .io_data_2_in_valid(PE_105_io_data_2_in_valid),
    .io_data_2_in_bits(PE_105_io_data_2_in_bits),
    .io_data_2_out_valid(PE_105_io_data_2_out_valid),
    .io_data_2_out_bits(PE_105_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_105_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_105_io_data_2_in_ready),
    .io_data_2_out_ready(PE_105_io_data_2_out_ready),
    .io_data_1_in_valid(PE_105_io_data_1_in_valid),
    .io_data_1_in_bits(PE_105_io_data_1_in_bits),
    .io_data_1_out_valid(PE_105_io_data_1_out_valid),
    .io_data_1_out_bits(PE_105_io_data_1_out_bits),
    .io_data_0_in_valid(PE_105_io_data_0_in_valid),
    .io_data_0_in_bits(PE_105_io_data_0_in_bits),
    .io_data_0_out_valid(PE_105_io_data_0_out_valid),
    .io_data_0_out_bits(PE_105_io_data_0_out_bits)
  );
  PE PE_106 ( // @[pe.scala 184:13]
    .clock(PE_106_clock),
    .reset(PE_106_reset),
    .io_data_2_in_valid(PE_106_io_data_2_in_valid),
    .io_data_2_in_bits(PE_106_io_data_2_in_bits),
    .io_data_2_out_valid(PE_106_io_data_2_out_valid),
    .io_data_2_out_bits(PE_106_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_106_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_106_io_data_2_in_ready),
    .io_data_2_out_ready(PE_106_io_data_2_out_ready),
    .io_data_1_in_valid(PE_106_io_data_1_in_valid),
    .io_data_1_in_bits(PE_106_io_data_1_in_bits),
    .io_data_1_out_valid(PE_106_io_data_1_out_valid),
    .io_data_1_out_bits(PE_106_io_data_1_out_bits),
    .io_data_0_in_valid(PE_106_io_data_0_in_valid),
    .io_data_0_in_bits(PE_106_io_data_0_in_bits),
    .io_data_0_out_valid(PE_106_io_data_0_out_valid),
    .io_data_0_out_bits(PE_106_io_data_0_out_bits)
  );
  PE PE_107 ( // @[pe.scala 184:13]
    .clock(PE_107_clock),
    .reset(PE_107_reset),
    .io_data_2_in_valid(PE_107_io_data_2_in_valid),
    .io_data_2_in_bits(PE_107_io_data_2_in_bits),
    .io_data_2_out_valid(PE_107_io_data_2_out_valid),
    .io_data_2_out_bits(PE_107_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_107_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_107_io_data_2_in_ready),
    .io_data_2_out_ready(PE_107_io_data_2_out_ready),
    .io_data_1_in_valid(PE_107_io_data_1_in_valid),
    .io_data_1_in_bits(PE_107_io_data_1_in_bits),
    .io_data_1_out_valid(PE_107_io_data_1_out_valid),
    .io_data_1_out_bits(PE_107_io_data_1_out_bits),
    .io_data_0_in_valid(PE_107_io_data_0_in_valid),
    .io_data_0_in_bits(PE_107_io_data_0_in_bits),
    .io_data_0_out_valid(PE_107_io_data_0_out_valid),
    .io_data_0_out_bits(PE_107_io_data_0_out_bits)
  );
  PE PE_108 ( // @[pe.scala 184:13]
    .clock(PE_108_clock),
    .reset(PE_108_reset),
    .io_data_2_in_valid(PE_108_io_data_2_in_valid),
    .io_data_2_in_bits(PE_108_io_data_2_in_bits),
    .io_data_2_out_valid(PE_108_io_data_2_out_valid),
    .io_data_2_out_bits(PE_108_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_108_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_108_io_data_2_in_ready),
    .io_data_2_out_ready(PE_108_io_data_2_out_ready),
    .io_data_1_in_valid(PE_108_io_data_1_in_valid),
    .io_data_1_in_bits(PE_108_io_data_1_in_bits),
    .io_data_1_out_valid(PE_108_io_data_1_out_valid),
    .io_data_1_out_bits(PE_108_io_data_1_out_bits),
    .io_data_0_in_valid(PE_108_io_data_0_in_valid),
    .io_data_0_in_bits(PE_108_io_data_0_in_bits),
    .io_data_0_out_valid(PE_108_io_data_0_out_valid),
    .io_data_0_out_bits(PE_108_io_data_0_out_bits)
  );
  PE PE_109 ( // @[pe.scala 184:13]
    .clock(PE_109_clock),
    .reset(PE_109_reset),
    .io_data_2_in_valid(PE_109_io_data_2_in_valid),
    .io_data_2_in_bits(PE_109_io_data_2_in_bits),
    .io_data_2_out_valid(PE_109_io_data_2_out_valid),
    .io_data_2_out_bits(PE_109_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_109_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_109_io_data_2_in_ready),
    .io_data_2_out_ready(PE_109_io_data_2_out_ready),
    .io_data_1_in_valid(PE_109_io_data_1_in_valid),
    .io_data_1_in_bits(PE_109_io_data_1_in_bits),
    .io_data_1_out_valid(PE_109_io_data_1_out_valid),
    .io_data_1_out_bits(PE_109_io_data_1_out_bits),
    .io_data_0_in_valid(PE_109_io_data_0_in_valid),
    .io_data_0_in_bits(PE_109_io_data_0_in_bits),
    .io_data_0_out_valid(PE_109_io_data_0_out_valid),
    .io_data_0_out_bits(PE_109_io_data_0_out_bits)
  );
  PE PE_110 ( // @[pe.scala 184:13]
    .clock(PE_110_clock),
    .reset(PE_110_reset),
    .io_data_2_in_valid(PE_110_io_data_2_in_valid),
    .io_data_2_in_bits(PE_110_io_data_2_in_bits),
    .io_data_2_out_valid(PE_110_io_data_2_out_valid),
    .io_data_2_out_bits(PE_110_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_110_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_110_io_data_2_in_ready),
    .io_data_2_out_ready(PE_110_io_data_2_out_ready),
    .io_data_1_in_valid(PE_110_io_data_1_in_valid),
    .io_data_1_in_bits(PE_110_io_data_1_in_bits),
    .io_data_1_out_valid(PE_110_io_data_1_out_valid),
    .io_data_1_out_bits(PE_110_io_data_1_out_bits),
    .io_data_0_in_valid(PE_110_io_data_0_in_valid),
    .io_data_0_in_bits(PE_110_io_data_0_in_bits),
    .io_data_0_out_valid(PE_110_io_data_0_out_valid),
    .io_data_0_out_bits(PE_110_io_data_0_out_bits)
  );
  PE PE_111 ( // @[pe.scala 184:13]
    .clock(PE_111_clock),
    .reset(PE_111_reset),
    .io_data_2_in_valid(PE_111_io_data_2_in_valid),
    .io_data_2_in_bits(PE_111_io_data_2_in_bits),
    .io_data_2_out_valid(PE_111_io_data_2_out_valid),
    .io_data_2_out_bits(PE_111_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_111_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_111_io_data_2_in_ready),
    .io_data_2_out_ready(PE_111_io_data_2_out_ready),
    .io_data_1_in_valid(PE_111_io_data_1_in_valid),
    .io_data_1_in_bits(PE_111_io_data_1_in_bits),
    .io_data_1_out_valid(PE_111_io_data_1_out_valid),
    .io_data_1_out_bits(PE_111_io_data_1_out_bits),
    .io_data_0_in_valid(PE_111_io_data_0_in_valid),
    .io_data_0_in_bits(PE_111_io_data_0_in_bits),
    .io_data_0_out_valid(PE_111_io_data_0_out_valid),
    .io_data_0_out_bits(PE_111_io_data_0_out_bits)
  );
  PE PE_112 ( // @[pe.scala 184:13]
    .clock(PE_112_clock),
    .reset(PE_112_reset),
    .io_data_2_in_valid(PE_112_io_data_2_in_valid),
    .io_data_2_in_bits(PE_112_io_data_2_in_bits),
    .io_data_2_out_valid(PE_112_io_data_2_out_valid),
    .io_data_2_out_bits(PE_112_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_112_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_112_io_data_2_in_ready),
    .io_data_2_out_ready(PE_112_io_data_2_out_ready),
    .io_data_1_in_valid(PE_112_io_data_1_in_valid),
    .io_data_1_in_bits(PE_112_io_data_1_in_bits),
    .io_data_1_out_valid(PE_112_io_data_1_out_valid),
    .io_data_1_out_bits(PE_112_io_data_1_out_bits),
    .io_data_0_in_valid(PE_112_io_data_0_in_valid),
    .io_data_0_in_bits(PE_112_io_data_0_in_bits),
    .io_data_0_out_valid(PE_112_io_data_0_out_valid),
    .io_data_0_out_bits(PE_112_io_data_0_out_bits)
  );
  PE PE_113 ( // @[pe.scala 184:13]
    .clock(PE_113_clock),
    .reset(PE_113_reset),
    .io_data_2_in_valid(PE_113_io_data_2_in_valid),
    .io_data_2_in_bits(PE_113_io_data_2_in_bits),
    .io_data_2_out_valid(PE_113_io_data_2_out_valid),
    .io_data_2_out_bits(PE_113_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_113_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_113_io_data_2_in_ready),
    .io_data_2_out_ready(PE_113_io_data_2_out_ready),
    .io_data_1_in_valid(PE_113_io_data_1_in_valid),
    .io_data_1_in_bits(PE_113_io_data_1_in_bits),
    .io_data_1_out_valid(PE_113_io_data_1_out_valid),
    .io_data_1_out_bits(PE_113_io_data_1_out_bits),
    .io_data_0_in_valid(PE_113_io_data_0_in_valid),
    .io_data_0_in_bits(PE_113_io_data_0_in_bits),
    .io_data_0_out_valid(PE_113_io_data_0_out_valid),
    .io_data_0_out_bits(PE_113_io_data_0_out_bits)
  );
  PE PE_114 ( // @[pe.scala 184:13]
    .clock(PE_114_clock),
    .reset(PE_114_reset),
    .io_data_2_in_valid(PE_114_io_data_2_in_valid),
    .io_data_2_in_bits(PE_114_io_data_2_in_bits),
    .io_data_2_out_valid(PE_114_io_data_2_out_valid),
    .io_data_2_out_bits(PE_114_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_114_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_114_io_data_2_in_ready),
    .io_data_2_out_ready(PE_114_io_data_2_out_ready),
    .io_data_1_in_valid(PE_114_io_data_1_in_valid),
    .io_data_1_in_bits(PE_114_io_data_1_in_bits),
    .io_data_1_out_valid(PE_114_io_data_1_out_valid),
    .io_data_1_out_bits(PE_114_io_data_1_out_bits),
    .io_data_0_in_valid(PE_114_io_data_0_in_valid),
    .io_data_0_in_bits(PE_114_io_data_0_in_bits),
    .io_data_0_out_valid(PE_114_io_data_0_out_valid),
    .io_data_0_out_bits(PE_114_io_data_0_out_bits)
  );
  PE PE_115 ( // @[pe.scala 184:13]
    .clock(PE_115_clock),
    .reset(PE_115_reset),
    .io_data_2_in_valid(PE_115_io_data_2_in_valid),
    .io_data_2_in_bits(PE_115_io_data_2_in_bits),
    .io_data_2_out_valid(PE_115_io_data_2_out_valid),
    .io_data_2_out_bits(PE_115_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_115_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_115_io_data_2_in_ready),
    .io_data_2_out_ready(PE_115_io_data_2_out_ready),
    .io_data_1_in_valid(PE_115_io_data_1_in_valid),
    .io_data_1_in_bits(PE_115_io_data_1_in_bits),
    .io_data_1_out_valid(PE_115_io_data_1_out_valid),
    .io_data_1_out_bits(PE_115_io_data_1_out_bits),
    .io_data_0_in_valid(PE_115_io_data_0_in_valid),
    .io_data_0_in_bits(PE_115_io_data_0_in_bits),
    .io_data_0_out_valid(PE_115_io_data_0_out_valid),
    .io_data_0_out_bits(PE_115_io_data_0_out_bits)
  );
  PE PE_116 ( // @[pe.scala 184:13]
    .clock(PE_116_clock),
    .reset(PE_116_reset),
    .io_data_2_in_valid(PE_116_io_data_2_in_valid),
    .io_data_2_in_bits(PE_116_io_data_2_in_bits),
    .io_data_2_out_valid(PE_116_io_data_2_out_valid),
    .io_data_2_out_bits(PE_116_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_116_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_116_io_data_2_in_ready),
    .io_data_2_out_ready(PE_116_io_data_2_out_ready),
    .io_data_1_in_valid(PE_116_io_data_1_in_valid),
    .io_data_1_in_bits(PE_116_io_data_1_in_bits),
    .io_data_1_out_valid(PE_116_io_data_1_out_valid),
    .io_data_1_out_bits(PE_116_io_data_1_out_bits),
    .io_data_0_in_valid(PE_116_io_data_0_in_valid),
    .io_data_0_in_bits(PE_116_io_data_0_in_bits),
    .io_data_0_out_valid(PE_116_io_data_0_out_valid),
    .io_data_0_out_bits(PE_116_io_data_0_out_bits)
  );
  PE PE_117 ( // @[pe.scala 184:13]
    .clock(PE_117_clock),
    .reset(PE_117_reset),
    .io_data_2_in_valid(PE_117_io_data_2_in_valid),
    .io_data_2_in_bits(PE_117_io_data_2_in_bits),
    .io_data_2_out_valid(PE_117_io_data_2_out_valid),
    .io_data_2_out_bits(PE_117_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_117_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_117_io_data_2_in_ready),
    .io_data_2_out_ready(PE_117_io_data_2_out_ready),
    .io_data_1_in_valid(PE_117_io_data_1_in_valid),
    .io_data_1_in_bits(PE_117_io_data_1_in_bits),
    .io_data_1_out_valid(PE_117_io_data_1_out_valid),
    .io_data_1_out_bits(PE_117_io_data_1_out_bits),
    .io_data_0_in_valid(PE_117_io_data_0_in_valid),
    .io_data_0_in_bits(PE_117_io_data_0_in_bits),
    .io_data_0_out_valid(PE_117_io_data_0_out_valid),
    .io_data_0_out_bits(PE_117_io_data_0_out_bits)
  );
  PE PE_118 ( // @[pe.scala 184:13]
    .clock(PE_118_clock),
    .reset(PE_118_reset),
    .io_data_2_in_valid(PE_118_io_data_2_in_valid),
    .io_data_2_in_bits(PE_118_io_data_2_in_bits),
    .io_data_2_out_valid(PE_118_io_data_2_out_valid),
    .io_data_2_out_bits(PE_118_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_118_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_118_io_data_2_in_ready),
    .io_data_2_out_ready(PE_118_io_data_2_out_ready),
    .io_data_1_in_valid(PE_118_io_data_1_in_valid),
    .io_data_1_in_bits(PE_118_io_data_1_in_bits),
    .io_data_1_out_valid(PE_118_io_data_1_out_valid),
    .io_data_1_out_bits(PE_118_io_data_1_out_bits),
    .io_data_0_in_valid(PE_118_io_data_0_in_valid),
    .io_data_0_in_bits(PE_118_io_data_0_in_bits),
    .io_data_0_out_valid(PE_118_io_data_0_out_valid),
    .io_data_0_out_bits(PE_118_io_data_0_out_bits)
  );
  PE PE_119 ( // @[pe.scala 184:13]
    .clock(PE_119_clock),
    .reset(PE_119_reset),
    .io_data_2_in_valid(PE_119_io_data_2_in_valid),
    .io_data_2_in_bits(PE_119_io_data_2_in_bits),
    .io_data_2_out_valid(PE_119_io_data_2_out_valid),
    .io_data_2_out_bits(PE_119_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_119_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_119_io_data_2_in_ready),
    .io_data_2_out_ready(PE_119_io_data_2_out_ready),
    .io_data_1_in_valid(PE_119_io_data_1_in_valid),
    .io_data_1_in_bits(PE_119_io_data_1_in_bits),
    .io_data_1_out_valid(PE_119_io_data_1_out_valid),
    .io_data_1_out_bits(PE_119_io_data_1_out_bits),
    .io_data_0_in_valid(PE_119_io_data_0_in_valid),
    .io_data_0_in_bits(PE_119_io_data_0_in_bits),
    .io_data_0_out_valid(PE_119_io_data_0_out_valid),
    .io_data_0_out_bits(PE_119_io_data_0_out_bits)
  );
  PE PE_120 ( // @[pe.scala 184:13]
    .clock(PE_120_clock),
    .reset(PE_120_reset),
    .io_data_2_in_valid(PE_120_io_data_2_in_valid),
    .io_data_2_in_bits(PE_120_io_data_2_in_bits),
    .io_data_2_out_valid(PE_120_io_data_2_out_valid),
    .io_data_2_out_bits(PE_120_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_120_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_120_io_data_2_in_ready),
    .io_data_2_out_ready(PE_120_io_data_2_out_ready),
    .io_data_1_in_valid(PE_120_io_data_1_in_valid),
    .io_data_1_in_bits(PE_120_io_data_1_in_bits),
    .io_data_1_out_valid(PE_120_io_data_1_out_valid),
    .io_data_1_out_bits(PE_120_io_data_1_out_bits),
    .io_data_0_in_valid(PE_120_io_data_0_in_valid),
    .io_data_0_in_bits(PE_120_io_data_0_in_bits),
    .io_data_0_out_valid(PE_120_io_data_0_out_valid),
    .io_data_0_out_bits(PE_120_io_data_0_out_bits)
  );
  PE PE_121 ( // @[pe.scala 184:13]
    .clock(PE_121_clock),
    .reset(PE_121_reset),
    .io_data_2_in_valid(PE_121_io_data_2_in_valid),
    .io_data_2_in_bits(PE_121_io_data_2_in_bits),
    .io_data_2_out_valid(PE_121_io_data_2_out_valid),
    .io_data_2_out_bits(PE_121_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_121_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_121_io_data_2_in_ready),
    .io_data_2_out_ready(PE_121_io_data_2_out_ready),
    .io_data_1_in_valid(PE_121_io_data_1_in_valid),
    .io_data_1_in_bits(PE_121_io_data_1_in_bits),
    .io_data_1_out_valid(PE_121_io_data_1_out_valid),
    .io_data_1_out_bits(PE_121_io_data_1_out_bits),
    .io_data_0_in_valid(PE_121_io_data_0_in_valid),
    .io_data_0_in_bits(PE_121_io_data_0_in_bits),
    .io_data_0_out_valid(PE_121_io_data_0_out_valid),
    .io_data_0_out_bits(PE_121_io_data_0_out_bits)
  );
  PE PE_122 ( // @[pe.scala 184:13]
    .clock(PE_122_clock),
    .reset(PE_122_reset),
    .io_data_2_in_valid(PE_122_io_data_2_in_valid),
    .io_data_2_in_bits(PE_122_io_data_2_in_bits),
    .io_data_2_out_valid(PE_122_io_data_2_out_valid),
    .io_data_2_out_bits(PE_122_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_122_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_122_io_data_2_in_ready),
    .io_data_2_out_ready(PE_122_io_data_2_out_ready),
    .io_data_1_in_valid(PE_122_io_data_1_in_valid),
    .io_data_1_in_bits(PE_122_io_data_1_in_bits),
    .io_data_1_out_valid(PE_122_io_data_1_out_valid),
    .io_data_1_out_bits(PE_122_io_data_1_out_bits),
    .io_data_0_in_valid(PE_122_io_data_0_in_valid),
    .io_data_0_in_bits(PE_122_io_data_0_in_bits),
    .io_data_0_out_valid(PE_122_io_data_0_out_valid),
    .io_data_0_out_bits(PE_122_io_data_0_out_bits)
  );
  PE PE_123 ( // @[pe.scala 184:13]
    .clock(PE_123_clock),
    .reset(PE_123_reset),
    .io_data_2_in_valid(PE_123_io_data_2_in_valid),
    .io_data_2_in_bits(PE_123_io_data_2_in_bits),
    .io_data_2_out_valid(PE_123_io_data_2_out_valid),
    .io_data_2_out_bits(PE_123_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_123_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_123_io_data_2_in_ready),
    .io_data_2_out_ready(PE_123_io_data_2_out_ready),
    .io_data_1_in_valid(PE_123_io_data_1_in_valid),
    .io_data_1_in_bits(PE_123_io_data_1_in_bits),
    .io_data_1_out_valid(PE_123_io_data_1_out_valid),
    .io_data_1_out_bits(PE_123_io_data_1_out_bits),
    .io_data_0_in_valid(PE_123_io_data_0_in_valid),
    .io_data_0_in_bits(PE_123_io_data_0_in_bits),
    .io_data_0_out_valid(PE_123_io_data_0_out_valid),
    .io_data_0_out_bits(PE_123_io_data_0_out_bits)
  );
  PE PE_124 ( // @[pe.scala 184:13]
    .clock(PE_124_clock),
    .reset(PE_124_reset),
    .io_data_2_in_valid(PE_124_io_data_2_in_valid),
    .io_data_2_in_bits(PE_124_io_data_2_in_bits),
    .io_data_2_out_valid(PE_124_io_data_2_out_valid),
    .io_data_2_out_bits(PE_124_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_124_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_124_io_data_2_in_ready),
    .io_data_2_out_ready(PE_124_io_data_2_out_ready),
    .io_data_1_in_valid(PE_124_io_data_1_in_valid),
    .io_data_1_in_bits(PE_124_io_data_1_in_bits),
    .io_data_1_out_valid(PE_124_io_data_1_out_valid),
    .io_data_1_out_bits(PE_124_io_data_1_out_bits),
    .io_data_0_in_valid(PE_124_io_data_0_in_valid),
    .io_data_0_in_bits(PE_124_io_data_0_in_bits),
    .io_data_0_out_valid(PE_124_io_data_0_out_valid),
    .io_data_0_out_bits(PE_124_io_data_0_out_bits)
  );
  PE PE_125 ( // @[pe.scala 184:13]
    .clock(PE_125_clock),
    .reset(PE_125_reset),
    .io_data_2_in_valid(PE_125_io_data_2_in_valid),
    .io_data_2_in_bits(PE_125_io_data_2_in_bits),
    .io_data_2_out_valid(PE_125_io_data_2_out_valid),
    .io_data_2_out_bits(PE_125_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_125_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_125_io_data_2_in_ready),
    .io_data_2_out_ready(PE_125_io_data_2_out_ready),
    .io_data_1_in_valid(PE_125_io_data_1_in_valid),
    .io_data_1_in_bits(PE_125_io_data_1_in_bits),
    .io_data_1_out_valid(PE_125_io_data_1_out_valid),
    .io_data_1_out_bits(PE_125_io_data_1_out_bits),
    .io_data_0_in_valid(PE_125_io_data_0_in_valid),
    .io_data_0_in_bits(PE_125_io_data_0_in_bits),
    .io_data_0_out_valid(PE_125_io_data_0_out_valid),
    .io_data_0_out_bits(PE_125_io_data_0_out_bits)
  );
  PE PE_126 ( // @[pe.scala 184:13]
    .clock(PE_126_clock),
    .reset(PE_126_reset),
    .io_data_2_in_valid(PE_126_io_data_2_in_valid),
    .io_data_2_in_bits(PE_126_io_data_2_in_bits),
    .io_data_2_out_valid(PE_126_io_data_2_out_valid),
    .io_data_2_out_bits(PE_126_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_126_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_126_io_data_2_in_ready),
    .io_data_2_out_ready(PE_126_io_data_2_out_ready),
    .io_data_1_in_valid(PE_126_io_data_1_in_valid),
    .io_data_1_in_bits(PE_126_io_data_1_in_bits),
    .io_data_1_out_valid(PE_126_io_data_1_out_valid),
    .io_data_1_out_bits(PE_126_io_data_1_out_bits),
    .io_data_0_in_valid(PE_126_io_data_0_in_valid),
    .io_data_0_in_bits(PE_126_io_data_0_in_bits),
    .io_data_0_out_valid(PE_126_io_data_0_out_valid),
    .io_data_0_out_bits(PE_126_io_data_0_out_bits)
  );
  PE PE_127 ( // @[pe.scala 184:13]
    .clock(PE_127_clock),
    .reset(PE_127_reset),
    .io_data_2_in_valid(PE_127_io_data_2_in_valid),
    .io_data_2_in_bits(PE_127_io_data_2_in_bits),
    .io_data_2_out_valid(PE_127_io_data_2_out_valid),
    .io_data_2_out_bits(PE_127_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_127_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_127_io_data_2_in_ready),
    .io_data_2_out_ready(PE_127_io_data_2_out_ready),
    .io_data_1_in_valid(PE_127_io_data_1_in_valid),
    .io_data_1_in_bits(PE_127_io_data_1_in_bits),
    .io_data_1_out_valid(PE_127_io_data_1_out_valid),
    .io_data_1_out_bits(PE_127_io_data_1_out_bits),
    .io_data_0_in_valid(PE_127_io_data_0_in_valid),
    .io_data_0_in_bits(PE_127_io_data_0_in_bits),
    .io_data_0_out_valid(PE_127_io_data_0_out_valid),
    .io_data_0_out_bits(PE_127_io_data_0_out_bits)
  );
  PE PE_128 ( // @[pe.scala 184:13]
    .clock(PE_128_clock),
    .reset(PE_128_reset),
    .io_data_2_in_valid(PE_128_io_data_2_in_valid),
    .io_data_2_in_bits(PE_128_io_data_2_in_bits),
    .io_data_2_out_valid(PE_128_io_data_2_out_valid),
    .io_data_2_out_bits(PE_128_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_128_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_128_io_data_2_in_ready),
    .io_data_2_out_ready(PE_128_io_data_2_out_ready),
    .io_data_1_in_valid(PE_128_io_data_1_in_valid),
    .io_data_1_in_bits(PE_128_io_data_1_in_bits),
    .io_data_1_out_valid(PE_128_io_data_1_out_valid),
    .io_data_1_out_bits(PE_128_io_data_1_out_bits),
    .io_data_0_in_valid(PE_128_io_data_0_in_valid),
    .io_data_0_in_bits(PE_128_io_data_0_in_bits),
    .io_data_0_out_valid(PE_128_io_data_0_out_valid),
    .io_data_0_out_bits(PE_128_io_data_0_out_bits)
  );
  PE PE_129 ( // @[pe.scala 184:13]
    .clock(PE_129_clock),
    .reset(PE_129_reset),
    .io_data_2_in_valid(PE_129_io_data_2_in_valid),
    .io_data_2_in_bits(PE_129_io_data_2_in_bits),
    .io_data_2_out_valid(PE_129_io_data_2_out_valid),
    .io_data_2_out_bits(PE_129_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_129_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_129_io_data_2_in_ready),
    .io_data_2_out_ready(PE_129_io_data_2_out_ready),
    .io_data_1_in_valid(PE_129_io_data_1_in_valid),
    .io_data_1_in_bits(PE_129_io_data_1_in_bits),
    .io_data_1_out_valid(PE_129_io_data_1_out_valid),
    .io_data_1_out_bits(PE_129_io_data_1_out_bits),
    .io_data_0_in_valid(PE_129_io_data_0_in_valid),
    .io_data_0_in_bits(PE_129_io_data_0_in_bits),
    .io_data_0_out_valid(PE_129_io_data_0_out_valid),
    .io_data_0_out_bits(PE_129_io_data_0_out_bits)
  );
  PE PE_130 ( // @[pe.scala 184:13]
    .clock(PE_130_clock),
    .reset(PE_130_reset),
    .io_data_2_in_valid(PE_130_io_data_2_in_valid),
    .io_data_2_in_bits(PE_130_io_data_2_in_bits),
    .io_data_2_out_valid(PE_130_io_data_2_out_valid),
    .io_data_2_out_bits(PE_130_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_130_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_130_io_data_2_in_ready),
    .io_data_2_out_ready(PE_130_io_data_2_out_ready),
    .io_data_1_in_valid(PE_130_io_data_1_in_valid),
    .io_data_1_in_bits(PE_130_io_data_1_in_bits),
    .io_data_1_out_valid(PE_130_io_data_1_out_valid),
    .io_data_1_out_bits(PE_130_io_data_1_out_bits),
    .io_data_0_in_valid(PE_130_io_data_0_in_valid),
    .io_data_0_in_bits(PE_130_io_data_0_in_bits),
    .io_data_0_out_valid(PE_130_io_data_0_out_valid),
    .io_data_0_out_bits(PE_130_io_data_0_out_bits)
  );
  PE PE_131 ( // @[pe.scala 184:13]
    .clock(PE_131_clock),
    .reset(PE_131_reset),
    .io_data_2_in_valid(PE_131_io_data_2_in_valid),
    .io_data_2_in_bits(PE_131_io_data_2_in_bits),
    .io_data_2_out_valid(PE_131_io_data_2_out_valid),
    .io_data_2_out_bits(PE_131_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_131_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_131_io_data_2_in_ready),
    .io_data_2_out_ready(PE_131_io_data_2_out_ready),
    .io_data_1_in_valid(PE_131_io_data_1_in_valid),
    .io_data_1_in_bits(PE_131_io_data_1_in_bits),
    .io_data_1_out_valid(PE_131_io_data_1_out_valid),
    .io_data_1_out_bits(PE_131_io_data_1_out_bits),
    .io_data_0_in_valid(PE_131_io_data_0_in_valid),
    .io_data_0_in_bits(PE_131_io_data_0_in_bits),
    .io_data_0_out_valid(PE_131_io_data_0_out_valid),
    .io_data_0_out_bits(PE_131_io_data_0_out_bits)
  );
  PE PE_132 ( // @[pe.scala 184:13]
    .clock(PE_132_clock),
    .reset(PE_132_reset),
    .io_data_2_in_valid(PE_132_io_data_2_in_valid),
    .io_data_2_in_bits(PE_132_io_data_2_in_bits),
    .io_data_2_out_valid(PE_132_io_data_2_out_valid),
    .io_data_2_out_bits(PE_132_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_132_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_132_io_data_2_in_ready),
    .io_data_2_out_ready(PE_132_io_data_2_out_ready),
    .io_data_1_in_valid(PE_132_io_data_1_in_valid),
    .io_data_1_in_bits(PE_132_io_data_1_in_bits),
    .io_data_1_out_valid(PE_132_io_data_1_out_valid),
    .io_data_1_out_bits(PE_132_io_data_1_out_bits),
    .io_data_0_in_valid(PE_132_io_data_0_in_valid),
    .io_data_0_in_bits(PE_132_io_data_0_in_bits),
    .io_data_0_out_valid(PE_132_io_data_0_out_valid),
    .io_data_0_out_bits(PE_132_io_data_0_out_bits)
  );
  PE PE_133 ( // @[pe.scala 184:13]
    .clock(PE_133_clock),
    .reset(PE_133_reset),
    .io_data_2_in_valid(PE_133_io_data_2_in_valid),
    .io_data_2_in_bits(PE_133_io_data_2_in_bits),
    .io_data_2_out_valid(PE_133_io_data_2_out_valid),
    .io_data_2_out_bits(PE_133_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_133_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_133_io_data_2_in_ready),
    .io_data_2_out_ready(PE_133_io_data_2_out_ready),
    .io_data_1_in_valid(PE_133_io_data_1_in_valid),
    .io_data_1_in_bits(PE_133_io_data_1_in_bits),
    .io_data_1_out_valid(PE_133_io_data_1_out_valid),
    .io_data_1_out_bits(PE_133_io_data_1_out_bits),
    .io_data_0_in_valid(PE_133_io_data_0_in_valid),
    .io_data_0_in_bits(PE_133_io_data_0_in_bits),
    .io_data_0_out_valid(PE_133_io_data_0_out_valid),
    .io_data_0_out_bits(PE_133_io_data_0_out_bits)
  );
  PE PE_134 ( // @[pe.scala 184:13]
    .clock(PE_134_clock),
    .reset(PE_134_reset),
    .io_data_2_in_valid(PE_134_io_data_2_in_valid),
    .io_data_2_in_bits(PE_134_io_data_2_in_bits),
    .io_data_2_out_valid(PE_134_io_data_2_out_valid),
    .io_data_2_out_bits(PE_134_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_134_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_134_io_data_2_in_ready),
    .io_data_2_out_ready(PE_134_io_data_2_out_ready),
    .io_data_1_in_valid(PE_134_io_data_1_in_valid),
    .io_data_1_in_bits(PE_134_io_data_1_in_bits),
    .io_data_1_out_valid(PE_134_io_data_1_out_valid),
    .io_data_1_out_bits(PE_134_io_data_1_out_bits),
    .io_data_0_in_valid(PE_134_io_data_0_in_valid),
    .io_data_0_in_bits(PE_134_io_data_0_in_bits),
    .io_data_0_out_valid(PE_134_io_data_0_out_valid),
    .io_data_0_out_bits(PE_134_io_data_0_out_bits)
  );
  PE PE_135 ( // @[pe.scala 184:13]
    .clock(PE_135_clock),
    .reset(PE_135_reset),
    .io_data_2_in_valid(PE_135_io_data_2_in_valid),
    .io_data_2_in_bits(PE_135_io_data_2_in_bits),
    .io_data_2_out_valid(PE_135_io_data_2_out_valid),
    .io_data_2_out_bits(PE_135_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_135_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_135_io_data_2_in_ready),
    .io_data_2_out_ready(PE_135_io_data_2_out_ready),
    .io_data_1_in_valid(PE_135_io_data_1_in_valid),
    .io_data_1_in_bits(PE_135_io_data_1_in_bits),
    .io_data_1_out_valid(PE_135_io_data_1_out_valid),
    .io_data_1_out_bits(PE_135_io_data_1_out_bits),
    .io_data_0_in_valid(PE_135_io_data_0_in_valid),
    .io_data_0_in_bits(PE_135_io_data_0_in_bits),
    .io_data_0_out_valid(PE_135_io_data_0_out_valid),
    .io_data_0_out_bits(PE_135_io_data_0_out_bits)
  );
  PE PE_136 ( // @[pe.scala 184:13]
    .clock(PE_136_clock),
    .reset(PE_136_reset),
    .io_data_2_in_valid(PE_136_io_data_2_in_valid),
    .io_data_2_in_bits(PE_136_io_data_2_in_bits),
    .io_data_2_out_valid(PE_136_io_data_2_out_valid),
    .io_data_2_out_bits(PE_136_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_136_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_136_io_data_2_in_ready),
    .io_data_2_out_ready(PE_136_io_data_2_out_ready),
    .io_data_1_in_valid(PE_136_io_data_1_in_valid),
    .io_data_1_in_bits(PE_136_io_data_1_in_bits),
    .io_data_1_out_valid(PE_136_io_data_1_out_valid),
    .io_data_1_out_bits(PE_136_io_data_1_out_bits),
    .io_data_0_in_valid(PE_136_io_data_0_in_valid),
    .io_data_0_in_bits(PE_136_io_data_0_in_bits),
    .io_data_0_out_valid(PE_136_io_data_0_out_valid),
    .io_data_0_out_bits(PE_136_io_data_0_out_bits)
  );
  PE PE_137 ( // @[pe.scala 184:13]
    .clock(PE_137_clock),
    .reset(PE_137_reset),
    .io_data_2_in_valid(PE_137_io_data_2_in_valid),
    .io_data_2_in_bits(PE_137_io_data_2_in_bits),
    .io_data_2_out_valid(PE_137_io_data_2_out_valid),
    .io_data_2_out_bits(PE_137_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_137_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_137_io_data_2_in_ready),
    .io_data_2_out_ready(PE_137_io_data_2_out_ready),
    .io_data_1_in_valid(PE_137_io_data_1_in_valid),
    .io_data_1_in_bits(PE_137_io_data_1_in_bits),
    .io_data_1_out_valid(PE_137_io_data_1_out_valid),
    .io_data_1_out_bits(PE_137_io_data_1_out_bits),
    .io_data_0_in_valid(PE_137_io_data_0_in_valid),
    .io_data_0_in_bits(PE_137_io_data_0_in_bits),
    .io_data_0_out_valid(PE_137_io_data_0_out_valid),
    .io_data_0_out_bits(PE_137_io_data_0_out_bits)
  );
  PE PE_138 ( // @[pe.scala 184:13]
    .clock(PE_138_clock),
    .reset(PE_138_reset),
    .io_data_2_in_valid(PE_138_io_data_2_in_valid),
    .io_data_2_in_bits(PE_138_io_data_2_in_bits),
    .io_data_2_out_valid(PE_138_io_data_2_out_valid),
    .io_data_2_out_bits(PE_138_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_138_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_138_io_data_2_in_ready),
    .io_data_2_out_ready(PE_138_io_data_2_out_ready),
    .io_data_1_in_valid(PE_138_io_data_1_in_valid),
    .io_data_1_in_bits(PE_138_io_data_1_in_bits),
    .io_data_1_out_valid(PE_138_io_data_1_out_valid),
    .io_data_1_out_bits(PE_138_io_data_1_out_bits),
    .io_data_0_in_valid(PE_138_io_data_0_in_valid),
    .io_data_0_in_bits(PE_138_io_data_0_in_bits),
    .io_data_0_out_valid(PE_138_io_data_0_out_valid),
    .io_data_0_out_bits(PE_138_io_data_0_out_bits)
  );
  PE PE_139 ( // @[pe.scala 184:13]
    .clock(PE_139_clock),
    .reset(PE_139_reset),
    .io_data_2_in_valid(PE_139_io_data_2_in_valid),
    .io_data_2_in_bits(PE_139_io_data_2_in_bits),
    .io_data_2_out_valid(PE_139_io_data_2_out_valid),
    .io_data_2_out_bits(PE_139_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_139_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_139_io_data_2_in_ready),
    .io_data_2_out_ready(PE_139_io_data_2_out_ready),
    .io_data_1_in_valid(PE_139_io_data_1_in_valid),
    .io_data_1_in_bits(PE_139_io_data_1_in_bits),
    .io_data_1_out_valid(PE_139_io_data_1_out_valid),
    .io_data_1_out_bits(PE_139_io_data_1_out_bits),
    .io_data_0_in_valid(PE_139_io_data_0_in_valid),
    .io_data_0_in_bits(PE_139_io_data_0_in_bits),
    .io_data_0_out_valid(PE_139_io_data_0_out_valid),
    .io_data_0_out_bits(PE_139_io_data_0_out_bits)
  );
  PE PE_140 ( // @[pe.scala 184:13]
    .clock(PE_140_clock),
    .reset(PE_140_reset),
    .io_data_2_in_valid(PE_140_io_data_2_in_valid),
    .io_data_2_in_bits(PE_140_io_data_2_in_bits),
    .io_data_2_out_valid(PE_140_io_data_2_out_valid),
    .io_data_2_out_bits(PE_140_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_140_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_140_io_data_2_in_ready),
    .io_data_2_out_ready(PE_140_io_data_2_out_ready),
    .io_data_1_in_valid(PE_140_io_data_1_in_valid),
    .io_data_1_in_bits(PE_140_io_data_1_in_bits),
    .io_data_1_out_valid(PE_140_io_data_1_out_valid),
    .io_data_1_out_bits(PE_140_io_data_1_out_bits),
    .io_data_0_in_valid(PE_140_io_data_0_in_valid),
    .io_data_0_in_bits(PE_140_io_data_0_in_bits),
    .io_data_0_out_valid(PE_140_io_data_0_out_valid),
    .io_data_0_out_bits(PE_140_io_data_0_out_bits)
  );
  PE PE_141 ( // @[pe.scala 184:13]
    .clock(PE_141_clock),
    .reset(PE_141_reset),
    .io_data_2_in_valid(PE_141_io_data_2_in_valid),
    .io_data_2_in_bits(PE_141_io_data_2_in_bits),
    .io_data_2_out_valid(PE_141_io_data_2_out_valid),
    .io_data_2_out_bits(PE_141_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_141_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_141_io_data_2_in_ready),
    .io_data_2_out_ready(PE_141_io_data_2_out_ready),
    .io_data_1_in_valid(PE_141_io_data_1_in_valid),
    .io_data_1_in_bits(PE_141_io_data_1_in_bits),
    .io_data_1_out_valid(PE_141_io_data_1_out_valid),
    .io_data_1_out_bits(PE_141_io_data_1_out_bits),
    .io_data_0_in_valid(PE_141_io_data_0_in_valid),
    .io_data_0_in_bits(PE_141_io_data_0_in_bits),
    .io_data_0_out_valid(PE_141_io_data_0_out_valid),
    .io_data_0_out_bits(PE_141_io_data_0_out_bits)
  );
  PE PE_142 ( // @[pe.scala 184:13]
    .clock(PE_142_clock),
    .reset(PE_142_reset),
    .io_data_2_in_valid(PE_142_io_data_2_in_valid),
    .io_data_2_in_bits(PE_142_io_data_2_in_bits),
    .io_data_2_out_valid(PE_142_io_data_2_out_valid),
    .io_data_2_out_bits(PE_142_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_142_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_142_io_data_2_in_ready),
    .io_data_2_out_ready(PE_142_io_data_2_out_ready),
    .io_data_1_in_valid(PE_142_io_data_1_in_valid),
    .io_data_1_in_bits(PE_142_io_data_1_in_bits),
    .io_data_1_out_valid(PE_142_io_data_1_out_valid),
    .io_data_1_out_bits(PE_142_io_data_1_out_bits),
    .io_data_0_in_valid(PE_142_io_data_0_in_valid),
    .io_data_0_in_bits(PE_142_io_data_0_in_bits),
    .io_data_0_out_valid(PE_142_io_data_0_out_valid),
    .io_data_0_out_bits(PE_142_io_data_0_out_bits)
  );
  PE PE_143 ( // @[pe.scala 184:13]
    .clock(PE_143_clock),
    .reset(PE_143_reset),
    .io_data_2_in_valid(PE_143_io_data_2_in_valid),
    .io_data_2_in_bits(PE_143_io_data_2_in_bits),
    .io_data_2_out_valid(PE_143_io_data_2_out_valid),
    .io_data_2_out_bits(PE_143_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_143_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_143_io_data_2_in_ready),
    .io_data_2_out_ready(PE_143_io_data_2_out_ready),
    .io_data_1_in_valid(PE_143_io_data_1_in_valid),
    .io_data_1_in_bits(PE_143_io_data_1_in_bits),
    .io_data_1_out_valid(PE_143_io_data_1_out_valid),
    .io_data_1_out_bits(PE_143_io_data_1_out_bits),
    .io_data_0_in_valid(PE_143_io_data_0_in_valid),
    .io_data_0_in_bits(PE_143_io_data_0_in_bits),
    .io_data_0_out_valid(PE_143_io_data_0_out_valid),
    .io_data_0_out_bits(PE_143_io_data_0_out_bits)
  );
  PE PE_144 ( // @[pe.scala 184:13]
    .clock(PE_144_clock),
    .reset(PE_144_reset),
    .io_data_2_in_valid(PE_144_io_data_2_in_valid),
    .io_data_2_in_bits(PE_144_io_data_2_in_bits),
    .io_data_2_out_valid(PE_144_io_data_2_out_valid),
    .io_data_2_out_bits(PE_144_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_144_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_144_io_data_2_in_ready),
    .io_data_2_out_ready(PE_144_io_data_2_out_ready),
    .io_data_1_in_valid(PE_144_io_data_1_in_valid),
    .io_data_1_in_bits(PE_144_io_data_1_in_bits),
    .io_data_1_out_valid(PE_144_io_data_1_out_valid),
    .io_data_1_out_bits(PE_144_io_data_1_out_bits),
    .io_data_0_in_valid(PE_144_io_data_0_in_valid),
    .io_data_0_in_bits(PE_144_io_data_0_in_bits),
    .io_data_0_out_valid(PE_144_io_data_0_out_valid),
    .io_data_0_out_bits(PE_144_io_data_0_out_bits)
  );
  PE PE_145 ( // @[pe.scala 184:13]
    .clock(PE_145_clock),
    .reset(PE_145_reset),
    .io_data_2_in_valid(PE_145_io_data_2_in_valid),
    .io_data_2_in_bits(PE_145_io_data_2_in_bits),
    .io_data_2_out_valid(PE_145_io_data_2_out_valid),
    .io_data_2_out_bits(PE_145_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_145_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_145_io_data_2_in_ready),
    .io_data_2_out_ready(PE_145_io_data_2_out_ready),
    .io_data_1_in_valid(PE_145_io_data_1_in_valid),
    .io_data_1_in_bits(PE_145_io_data_1_in_bits),
    .io_data_1_out_valid(PE_145_io_data_1_out_valid),
    .io_data_1_out_bits(PE_145_io_data_1_out_bits),
    .io_data_0_in_valid(PE_145_io_data_0_in_valid),
    .io_data_0_in_bits(PE_145_io_data_0_in_bits),
    .io_data_0_out_valid(PE_145_io_data_0_out_valid),
    .io_data_0_out_bits(PE_145_io_data_0_out_bits)
  );
  PE PE_146 ( // @[pe.scala 184:13]
    .clock(PE_146_clock),
    .reset(PE_146_reset),
    .io_data_2_in_valid(PE_146_io_data_2_in_valid),
    .io_data_2_in_bits(PE_146_io_data_2_in_bits),
    .io_data_2_out_valid(PE_146_io_data_2_out_valid),
    .io_data_2_out_bits(PE_146_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_146_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_146_io_data_2_in_ready),
    .io_data_2_out_ready(PE_146_io_data_2_out_ready),
    .io_data_1_in_valid(PE_146_io_data_1_in_valid),
    .io_data_1_in_bits(PE_146_io_data_1_in_bits),
    .io_data_1_out_valid(PE_146_io_data_1_out_valid),
    .io_data_1_out_bits(PE_146_io_data_1_out_bits),
    .io_data_0_in_valid(PE_146_io_data_0_in_valid),
    .io_data_0_in_bits(PE_146_io_data_0_in_bits),
    .io_data_0_out_valid(PE_146_io_data_0_out_valid),
    .io_data_0_out_bits(PE_146_io_data_0_out_bits)
  );
  PE PE_147 ( // @[pe.scala 184:13]
    .clock(PE_147_clock),
    .reset(PE_147_reset),
    .io_data_2_in_valid(PE_147_io_data_2_in_valid),
    .io_data_2_in_bits(PE_147_io_data_2_in_bits),
    .io_data_2_out_valid(PE_147_io_data_2_out_valid),
    .io_data_2_out_bits(PE_147_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_147_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_147_io_data_2_in_ready),
    .io_data_2_out_ready(PE_147_io_data_2_out_ready),
    .io_data_1_in_valid(PE_147_io_data_1_in_valid),
    .io_data_1_in_bits(PE_147_io_data_1_in_bits),
    .io_data_1_out_valid(PE_147_io_data_1_out_valid),
    .io_data_1_out_bits(PE_147_io_data_1_out_bits),
    .io_data_0_in_valid(PE_147_io_data_0_in_valid),
    .io_data_0_in_bits(PE_147_io_data_0_in_bits),
    .io_data_0_out_valid(PE_147_io_data_0_out_valid),
    .io_data_0_out_bits(PE_147_io_data_0_out_bits)
  );
  PE PE_148 ( // @[pe.scala 184:13]
    .clock(PE_148_clock),
    .reset(PE_148_reset),
    .io_data_2_in_valid(PE_148_io_data_2_in_valid),
    .io_data_2_in_bits(PE_148_io_data_2_in_bits),
    .io_data_2_out_valid(PE_148_io_data_2_out_valid),
    .io_data_2_out_bits(PE_148_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_148_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_148_io_data_2_in_ready),
    .io_data_2_out_ready(PE_148_io_data_2_out_ready),
    .io_data_1_in_valid(PE_148_io_data_1_in_valid),
    .io_data_1_in_bits(PE_148_io_data_1_in_bits),
    .io_data_1_out_valid(PE_148_io_data_1_out_valid),
    .io_data_1_out_bits(PE_148_io_data_1_out_bits),
    .io_data_0_in_valid(PE_148_io_data_0_in_valid),
    .io_data_0_in_bits(PE_148_io_data_0_in_bits),
    .io_data_0_out_valid(PE_148_io_data_0_out_valid),
    .io_data_0_out_bits(PE_148_io_data_0_out_bits)
  );
  PE PE_149 ( // @[pe.scala 184:13]
    .clock(PE_149_clock),
    .reset(PE_149_reset),
    .io_data_2_in_valid(PE_149_io_data_2_in_valid),
    .io_data_2_in_bits(PE_149_io_data_2_in_bits),
    .io_data_2_out_valid(PE_149_io_data_2_out_valid),
    .io_data_2_out_bits(PE_149_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_149_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_149_io_data_2_in_ready),
    .io_data_2_out_ready(PE_149_io_data_2_out_ready),
    .io_data_1_in_valid(PE_149_io_data_1_in_valid),
    .io_data_1_in_bits(PE_149_io_data_1_in_bits),
    .io_data_1_out_valid(PE_149_io_data_1_out_valid),
    .io_data_1_out_bits(PE_149_io_data_1_out_bits),
    .io_data_0_in_valid(PE_149_io_data_0_in_valid),
    .io_data_0_in_bits(PE_149_io_data_0_in_bits),
    .io_data_0_out_valid(PE_149_io_data_0_out_valid),
    .io_data_0_out_bits(PE_149_io_data_0_out_bits)
  );
  PE PE_150 ( // @[pe.scala 184:13]
    .clock(PE_150_clock),
    .reset(PE_150_reset),
    .io_data_2_in_valid(PE_150_io_data_2_in_valid),
    .io_data_2_in_bits(PE_150_io_data_2_in_bits),
    .io_data_2_out_valid(PE_150_io_data_2_out_valid),
    .io_data_2_out_bits(PE_150_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_150_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_150_io_data_2_in_ready),
    .io_data_2_out_ready(PE_150_io_data_2_out_ready),
    .io_data_1_in_valid(PE_150_io_data_1_in_valid),
    .io_data_1_in_bits(PE_150_io_data_1_in_bits),
    .io_data_1_out_valid(PE_150_io_data_1_out_valid),
    .io_data_1_out_bits(PE_150_io_data_1_out_bits),
    .io_data_0_in_valid(PE_150_io_data_0_in_valid),
    .io_data_0_in_bits(PE_150_io_data_0_in_bits),
    .io_data_0_out_valid(PE_150_io_data_0_out_valid),
    .io_data_0_out_bits(PE_150_io_data_0_out_bits)
  );
  PE PE_151 ( // @[pe.scala 184:13]
    .clock(PE_151_clock),
    .reset(PE_151_reset),
    .io_data_2_in_valid(PE_151_io_data_2_in_valid),
    .io_data_2_in_bits(PE_151_io_data_2_in_bits),
    .io_data_2_out_valid(PE_151_io_data_2_out_valid),
    .io_data_2_out_bits(PE_151_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_151_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_151_io_data_2_in_ready),
    .io_data_2_out_ready(PE_151_io_data_2_out_ready),
    .io_data_1_in_valid(PE_151_io_data_1_in_valid),
    .io_data_1_in_bits(PE_151_io_data_1_in_bits),
    .io_data_1_out_valid(PE_151_io_data_1_out_valid),
    .io_data_1_out_bits(PE_151_io_data_1_out_bits),
    .io_data_0_in_valid(PE_151_io_data_0_in_valid),
    .io_data_0_in_bits(PE_151_io_data_0_in_bits),
    .io_data_0_out_valid(PE_151_io_data_0_out_valid),
    .io_data_0_out_bits(PE_151_io_data_0_out_bits)
  );
  PE PE_152 ( // @[pe.scala 184:13]
    .clock(PE_152_clock),
    .reset(PE_152_reset),
    .io_data_2_in_valid(PE_152_io_data_2_in_valid),
    .io_data_2_in_bits(PE_152_io_data_2_in_bits),
    .io_data_2_out_valid(PE_152_io_data_2_out_valid),
    .io_data_2_out_bits(PE_152_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_152_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_152_io_data_2_in_ready),
    .io_data_2_out_ready(PE_152_io_data_2_out_ready),
    .io_data_1_in_valid(PE_152_io_data_1_in_valid),
    .io_data_1_in_bits(PE_152_io_data_1_in_bits),
    .io_data_1_out_valid(PE_152_io_data_1_out_valid),
    .io_data_1_out_bits(PE_152_io_data_1_out_bits),
    .io_data_0_in_valid(PE_152_io_data_0_in_valid),
    .io_data_0_in_bits(PE_152_io_data_0_in_bits),
    .io_data_0_out_valid(PE_152_io_data_0_out_valid),
    .io_data_0_out_bits(PE_152_io_data_0_out_bits)
  );
  PE PE_153 ( // @[pe.scala 184:13]
    .clock(PE_153_clock),
    .reset(PE_153_reset),
    .io_data_2_in_valid(PE_153_io_data_2_in_valid),
    .io_data_2_in_bits(PE_153_io_data_2_in_bits),
    .io_data_2_out_valid(PE_153_io_data_2_out_valid),
    .io_data_2_out_bits(PE_153_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_153_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_153_io_data_2_in_ready),
    .io_data_2_out_ready(PE_153_io_data_2_out_ready),
    .io_data_1_in_valid(PE_153_io_data_1_in_valid),
    .io_data_1_in_bits(PE_153_io_data_1_in_bits),
    .io_data_1_out_valid(PE_153_io_data_1_out_valid),
    .io_data_1_out_bits(PE_153_io_data_1_out_bits),
    .io_data_0_in_valid(PE_153_io_data_0_in_valid),
    .io_data_0_in_bits(PE_153_io_data_0_in_bits),
    .io_data_0_out_valid(PE_153_io_data_0_out_valid),
    .io_data_0_out_bits(PE_153_io_data_0_out_bits)
  );
  PE PE_154 ( // @[pe.scala 184:13]
    .clock(PE_154_clock),
    .reset(PE_154_reset),
    .io_data_2_in_valid(PE_154_io_data_2_in_valid),
    .io_data_2_in_bits(PE_154_io_data_2_in_bits),
    .io_data_2_out_valid(PE_154_io_data_2_out_valid),
    .io_data_2_out_bits(PE_154_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_154_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_154_io_data_2_in_ready),
    .io_data_2_out_ready(PE_154_io_data_2_out_ready),
    .io_data_1_in_valid(PE_154_io_data_1_in_valid),
    .io_data_1_in_bits(PE_154_io_data_1_in_bits),
    .io_data_1_out_valid(PE_154_io_data_1_out_valid),
    .io_data_1_out_bits(PE_154_io_data_1_out_bits),
    .io_data_0_in_valid(PE_154_io_data_0_in_valid),
    .io_data_0_in_bits(PE_154_io_data_0_in_bits),
    .io_data_0_out_valid(PE_154_io_data_0_out_valid),
    .io_data_0_out_bits(PE_154_io_data_0_out_bits)
  );
  PE PE_155 ( // @[pe.scala 184:13]
    .clock(PE_155_clock),
    .reset(PE_155_reset),
    .io_data_2_in_valid(PE_155_io_data_2_in_valid),
    .io_data_2_in_bits(PE_155_io_data_2_in_bits),
    .io_data_2_out_valid(PE_155_io_data_2_out_valid),
    .io_data_2_out_bits(PE_155_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_155_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_155_io_data_2_in_ready),
    .io_data_2_out_ready(PE_155_io_data_2_out_ready),
    .io_data_1_in_valid(PE_155_io_data_1_in_valid),
    .io_data_1_in_bits(PE_155_io_data_1_in_bits),
    .io_data_1_out_valid(PE_155_io_data_1_out_valid),
    .io_data_1_out_bits(PE_155_io_data_1_out_bits),
    .io_data_0_in_valid(PE_155_io_data_0_in_valid),
    .io_data_0_in_bits(PE_155_io_data_0_in_bits),
    .io_data_0_out_valid(PE_155_io_data_0_out_valid),
    .io_data_0_out_bits(PE_155_io_data_0_out_bits)
  );
  PE PE_156 ( // @[pe.scala 184:13]
    .clock(PE_156_clock),
    .reset(PE_156_reset),
    .io_data_2_in_valid(PE_156_io_data_2_in_valid),
    .io_data_2_in_bits(PE_156_io_data_2_in_bits),
    .io_data_2_out_valid(PE_156_io_data_2_out_valid),
    .io_data_2_out_bits(PE_156_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_156_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_156_io_data_2_in_ready),
    .io_data_2_out_ready(PE_156_io_data_2_out_ready),
    .io_data_1_in_valid(PE_156_io_data_1_in_valid),
    .io_data_1_in_bits(PE_156_io_data_1_in_bits),
    .io_data_1_out_valid(PE_156_io_data_1_out_valid),
    .io_data_1_out_bits(PE_156_io_data_1_out_bits),
    .io_data_0_in_valid(PE_156_io_data_0_in_valid),
    .io_data_0_in_bits(PE_156_io_data_0_in_bits),
    .io_data_0_out_valid(PE_156_io_data_0_out_valid),
    .io_data_0_out_bits(PE_156_io_data_0_out_bits)
  );
  PE PE_157 ( // @[pe.scala 184:13]
    .clock(PE_157_clock),
    .reset(PE_157_reset),
    .io_data_2_in_valid(PE_157_io_data_2_in_valid),
    .io_data_2_in_bits(PE_157_io_data_2_in_bits),
    .io_data_2_out_valid(PE_157_io_data_2_out_valid),
    .io_data_2_out_bits(PE_157_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_157_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_157_io_data_2_in_ready),
    .io_data_2_out_ready(PE_157_io_data_2_out_ready),
    .io_data_1_in_valid(PE_157_io_data_1_in_valid),
    .io_data_1_in_bits(PE_157_io_data_1_in_bits),
    .io_data_1_out_valid(PE_157_io_data_1_out_valid),
    .io_data_1_out_bits(PE_157_io_data_1_out_bits),
    .io_data_0_in_valid(PE_157_io_data_0_in_valid),
    .io_data_0_in_bits(PE_157_io_data_0_in_bits),
    .io_data_0_out_valid(PE_157_io_data_0_out_valid),
    .io_data_0_out_bits(PE_157_io_data_0_out_bits)
  );
  PE PE_158 ( // @[pe.scala 184:13]
    .clock(PE_158_clock),
    .reset(PE_158_reset),
    .io_data_2_in_valid(PE_158_io_data_2_in_valid),
    .io_data_2_in_bits(PE_158_io_data_2_in_bits),
    .io_data_2_out_valid(PE_158_io_data_2_out_valid),
    .io_data_2_out_bits(PE_158_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_158_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_158_io_data_2_in_ready),
    .io_data_2_out_ready(PE_158_io_data_2_out_ready),
    .io_data_1_in_valid(PE_158_io_data_1_in_valid),
    .io_data_1_in_bits(PE_158_io_data_1_in_bits),
    .io_data_1_out_valid(PE_158_io_data_1_out_valid),
    .io_data_1_out_bits(PE_158_io_data_1_out_bits),
    .io_data_0_in_valid(PE_158_io_data_0_in_valid),
    .io_data_0_in_bits(PE_158_io_data_0_in_bits),
    .io_data_0_out_valid(PE_158_io_data_0_out_valid),
    .io_data_0_out_bits(PE_158_io_data_0_out_bits)
  );
  PE PE_159 ( // @[pe.scala 184:13]
    .clock(PE_159_clock),
    .reset(PE_159_reset),
    .io_data_2_in_valid(PE_159_io_data_2_in_valid),
    .io_data_2_in_bits(PE_159_io_data_2_in_bits),
    .io_data_2_out_valid(PE_159_io_data_2_out_valid),
    .io_data_2_out_bits(PE_159_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_159_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_159_io_data_2_in_ready),
    .io_data_2_out_ready(PE_159_io_data_2_out_ready),
    .io_data_1_in_valid(PE_159_io_data_1_in_valid),
    .io_data_1_in_bits(PE_159_io_data_1_in_bits),
    .io_data_1_out_valid(PE_159_io_data_1_out_valid),
    .io_data_1_out_bits(PE_159_io_data_1_out_bits),
    .io_data_0_in_valid(PE_159_io_data_0_in_valid),
    .io_data_0_in_bits(PE_159_io_data_0_in_bits),
    .io_data_0_out_valid(PE_159_io_data_0_out_valid),
    .io_data_0_out_bits(PE_159_io_data_0_out_bits)
  );
  PE PE_160 ( // @[pe.scala 184:13]
    .clock(PE_160_clock),
    .reset(PE_160_reset),
    .io_data_2_in_valid(PE_160_io_data_2_in_valid),
    .io_data_2_in_bits(PE_160_io_data_2_in_bits),
    .io_data_2_out_valid(PE_160_io_data_2_out_valid),
    .io_data_2_out_bits(PE_160_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_160_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_160_io_data_2_in_ready),
    .io_data_2_out_ready(PE_160_io_data_2_out_ready),
    .io_data_1_in_valid(PE_160_io_data_1_in_valid),
    .io_data_1_in_bits(PE_160_io_data_1_in_bits),
    .io_data_1_out_valid(PE_160_io_data_1_out_valid),
    .io_data_1_out_bits(PE_160_io_data_1_out_bits),
    .io_data_0_in_valid(PE_160_io_data_0_in_valid),
    .io_data_0_in_bits(PE_160_io_data_0_in_bits),
    .io_data_0_out_valid(PE_160_io_data_0_out_valid),
    .io_data_0_out_bits(PE_160_io_data_0_out_bits)
  );
  PE PE_161 ( // @[pe.scala 184:13]
    .clock(PE_161_clock),
    .reset(PE_161_reset),
    .io_data_2_in_valid(PE_161_io_data_2_in_valid),
    .io_data_2_in_bits(PE_161_io_data_2_in_bits),
    .io_data_2_out_valid(PE_161_io_data_2_out_valid),
    .io_data_2_out_bits(PE_161_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_161_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_161_io_data_2_in_ready),
    .io_data_2_out_ready(PE_161_io_data_2_out_ready),
    .io_data_1_in_valid(PE_161_io_data_1_in_valid),
    .io_data_1_in_bits(PE_161_io_data_1_in_bits),
    .io_data_1_out_valid(PE_161_io_data_1_out_valid),
    .io_data_1_out_bits(PE_161_io_data_1_out_bits),
    .io_data_0_in_valid(PE_161_io_data_0_in_valid),
    .io_data_0_in_bits(PE_161_io_data_0_in_bits),
    .io_data_0_out_valid(PE_161_io_data_0_out_valid),
    .io_data_0_out_bits(PE_161_io_data_0_out_bits)
  );
  PE PE_162 ( // @[pe.scala 184:13]
    .clock(PE_162_clock),
    .reset(PE_162_reset),
    .io_data_2_in_valid(PE_162_io_data_2_in_valid),
    .io_data_2_in_bits(PE_162_io_data_2_in_bits),
    .io_data_2_out_valid(PE_162_io_data_2_out_valid),
    .io_data_2_out_bits(PE_162_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_162_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_162_io_data_2_in_ready),
    .io_data_2_out_ready(PE_162_io_data_2_out_ready),
    .io_data_1_in_valid(PE_162_io_data_1_in_valid),
    .io_data_1_in_bits(PE_162_io_data_1_in_bits),
    .io_data_1_out_valid(PE_162_io_data_1_out_valid),
    .io_data_1_out_bits(PE_162_io_data_1_out_bits),
    .io_data_0_in_valid(PE_162_io_data_0_in_valid),
    .io_data_0_in_bits(PE_162_io_data_0_in_bits),
    .io_data_0_out_valid(PE_162_io_data_0_out_valid),
    .io_data_0_out_bits(PE_162_io_data_0_out_bits)
  );
  PE PE_163 ( // @[pe.scala 184:13]
    .clock(PE_163_clock),
    .reset(PE_163_reset),
    .io_data_2_in_valid(PE_163_io_data_2_in_valid),
    .io_data_2_in_bits(PE_163_io_data_2_in_bits),
    .io_data_2_out_valid(PE_163_io_data_2_out_valid),
    .io_data_2_out_bits(PE_163_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_163_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_163_io_data_2_in_ready),
    .io_data_2_out_ready(PE_163_io_data_2_out_ready),
    .io_data_1_in_valid(PE_163_io_data_1_in_valid),
    .io_data_1_in_bits(PE_163_io_data_1_in_bits),
    .io_data_1_out_valid(PE_163_io_data_1_out_valid),
    .io_data_1_out_bits(PE_163_io_data_1_out_bits),
    .io_data_0_in_valid(PE_163_io_data_0_in_valid),
    .io_data_0_in_bits(PE_163_io_data_0_in_bits),
    .io_data_0_out_valid(PE_163_io_data_0_out_valid),
    .io_data_0_out_bits(PE_163_io_data_0_out_bits)
  );
  PE PE_164 ( // @[pe.scala 184:13]
    .clock(PE_164_clock),
    .reset(PE_164_reset),
    .io_data_2_in_valid(PE_164_io_data_2_in_valid),
    .io_data_2_in_bits(PE_164_io_data_2_in_bits),
    .io_data_2_out_valid(PE_164_io_data_2_out_valid),
    .io_data_2_out_bits(PE_164_io_data_2_out_bits),
    .io_data_2_sig_stat2trans(PE_164_io_data_2_sig_stat2trans),
    .io_data_2_in_ready(PE_164_io_data_2_in_ready),
    .io_data_2_out_ready(PE_164_io_data_2_out_ready),
    .io_data_1_in_valid(PE_164_io_data_1_in_valid),
    .io_data_1_in_bits(PE_164_io_data_1_in_bits),
    .io_data_1_out_valid(PE_164_io_data_1_out_valid),
    .io_data_1_out_bits(PE_164_io_data_1_out_bits),
    .io_data_0_in_valid(PE_164_io_data_0_in_valid),
    .io_data_0_in_bits(PE_164_io_data_0_in_bits),
    .io_data_0_out_valid(PE_164_io_data_0_out_valid),
    .io_data_0_out_bits(PE_164_io_data_0_out_bits)
  );
  PENetwork PENetwork ( // @[pe.scala 227:13]
    .io_to_pes_0_in_valid(PENetwork_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_io_to_pes_14_in_bits),
    .io_to_mem_valid(PENetwork_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_io_to_mem_bits)
  );
  PENetwork PENetwork_1 ( // @[pe.scala 227:13]
    .io_to_pes_0_in_valid(PENetwork_1_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_1_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_1_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_1_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_1_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_1_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_1_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_1_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_1_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_1_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_1_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_1_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_1_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_1_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_1_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_1_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_1_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_1_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_1_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_1_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_1_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_1_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_1_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_1_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_1_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_1_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_1_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_1_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_1_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_1_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_1_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_1_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_1_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_1_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_1_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_1_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_1_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_1_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_1_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_1_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_1_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_1_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_1_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_1_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_1_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_1_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_1_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_1_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_1_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_1_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_1_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_1_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_1_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_1_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_1_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_1_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_1_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_1_io_to_pes_14_in_bits),
    .io_to_mem_valid(PENetwork_1_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_1_io_to_mem_bits)
  );
  PENetwork PENetwork_2 ( // @[pe.scala 227:13]
    .io_to_pes_0_in_valid(PENetwork_2_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_2_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_2_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_2_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_2_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_2_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_2_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_2_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_2_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_2_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_2_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_2_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_2_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_2_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_2_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_2_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_2_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_2_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_2_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_2_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_2_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_2_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_2_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_2_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_2_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_2_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_2_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_2_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_2_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_2_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_2_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_2_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_2_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_2_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_2_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_2_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_2_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_2_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_2_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_2_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_2_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_2_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_2_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_2_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_2_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_2_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_2_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_2_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_2_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_2_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_2_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_2_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_2_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_2_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_2_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_2_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_2_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_2_io_to_pes_14_in_bits),
    .io_to_mem_valid(PENetwork_2_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_2_io_to_mem_bits)
  );
  PENetwork PENetwork_3 ( // @[pe.scala 227:13]
    .io_to_pes_0_in_valid(PENetwork_3_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_3_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_3_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_3_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_3_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_3_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_3_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_3_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_3_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_3_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_3_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_3_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_3_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_3_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_3_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_3_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_3_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_3_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_3_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_3_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_3_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_3_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_3_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_3_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_3_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_3_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_3_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_3_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_3_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_3_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_3_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_3_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_3_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_3_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_3_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_3_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_3_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_3_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_3_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_3_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_3_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_3_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_3_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_3_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_3_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_3_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_3_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_3_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_3_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_3_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_3_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_3_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_3_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_3_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_3_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_3_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_3_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_3_io_to_pes_14_in_bits),
    .io_to_mem_valid(PENetwork_3_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_3_io_to_mem_bits)
  );
  PENetwork PENetwork_4 ( // @[pe.scala 227:13]
    .io_to_pes_0_in_valid(PENetwork_4_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_4_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_4_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_4_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_4_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_4_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_4_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_4_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_4_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_4_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_4_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_4_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_4_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_4_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_4_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_4_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_4_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_4_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_4_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_4_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_4_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_4_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_4_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_4_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_4_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_4_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_4_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_4_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_4_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_4_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_4_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_4_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_4_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_4_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_4_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_4_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_4_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_4_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_4_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_4_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_4_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_4_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_4_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_4_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_4_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_4_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_4_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_4_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_4_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_4_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_4_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_4_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_4_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_4_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_4_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_4_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_4_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_4_io_to_pes_14_in_bits),
    .io_to_mem_valid(PENetwork_4_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_4_io_to_mem_bits)
  );
  PENetwork PENetwork_5 ( // @[pe.scala 227:13]
    .io_to_pes_0_in_valid(PENetwork_5_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_5_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_5_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_5_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_5_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_5_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_5_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_5_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_5_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_5_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_5_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_5_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_5_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_5_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_5_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_5_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_5_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_5_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_5_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_5_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_5_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_5_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_5_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_5_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_5_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_5_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_5_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_5_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_5_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_5_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_5_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_5_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_5_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_5_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_5_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_5_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_5_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_5_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_5_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_5_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_5_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_5_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_5_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_5_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_5_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_5_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_5_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_5_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_5_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_5_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_5_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_5_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_5_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_5_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_5_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_5_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_5_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_5_io_to_pes_14_in_bits),
    .io_to_mem_valid(PENetwork_5_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_5_io_to_mem_bits)
  );
  PENetwork PENetwork_6 ( // @[pe.scala 227:13]
    .io_to_pes_0_in_valid(PENetwork_6_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_6_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_6_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_6_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_6_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_6_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_6_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_6_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_6_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_6_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_6_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_6_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_6_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_6_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_6_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_6_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_6_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_6_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_6_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_6_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_6_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_6_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_6_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_6_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_6_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_6_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_6_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_6_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_6_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_6_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_6_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_6_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_6_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_6_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_6_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_6_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_6_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_6_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_6_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_6_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_6_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_6_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_6_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_6_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_6_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_6_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_6_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_6_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_6_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_6_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_6_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_6_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_6_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_6_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_6_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_6_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_6_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_6_io_to_pes_14_in_bits),
    .io_to_mem_valid(PENetwork_6_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_6_io_to_mem_bits)
  );
  PENetwork PENetwork_7 ( // @[pe.scala 227:13]
    .io_to_pes_0_in_valid(PENetwork_7_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_7_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_7_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_7_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_7_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_7_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_7_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_7_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_7_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_7_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_7_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_7_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_7_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_7_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_7_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_7_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_7_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_7_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_7_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_7_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_7_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_7_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_7_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_7_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_7_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_7_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_7_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_7_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_7_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_7_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_7_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_7_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_7_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_7_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_7_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_7_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_7_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_7_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_7_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_7_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_7_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_7_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_7_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_7_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_7_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_7_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_7_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_7_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_7_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_7_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_7_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_7_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_7_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_7_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_7_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_7_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_7_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_7_io_to_pes_14_in_bits),
    .io_to_mem_valid(PENetwork_7_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_7_io_to_mem_bits)
  );
  PENetwork PENetwork_8 ( // @[pe.scala 227:13]
    .io_to_pes_0_in_valid(PENetwork_8_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_8_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_8_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_8_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_8_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_8_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_8_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_8_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_8_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_8_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_8_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_8_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_8_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_8_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_8_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_8_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_8_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_8_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_8_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_8_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_8_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_8_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_8_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_8_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_8_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_8_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_8_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_8_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_8_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_8_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_8_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_8_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_8_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_8_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_8_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_8_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_8_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_8_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_8_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_8_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_8_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_8_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_8_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_8_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_8_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_8_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_8_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_8_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_8_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_8_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_8_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_8_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_8_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_8_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_8_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_8_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_8_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_8_io_to_pes_14_in_bits),
    .io_to_mem_valid(PENetwork_8_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_8_io_to_mem_bits)
  );
  PENetwork PENetwork_9 ( // @[pe.scala 227:13]
    .io_to_pes_0_in_valid(PENetwork_9_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_9_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_9_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_9_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_9_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_9_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_9_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_9_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_9_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_9_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_9_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_9_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_9_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_9_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_9_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_9_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_9_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_9_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_9_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_9_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_9_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_9_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_9_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_9_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_9_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_9_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_9_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_9_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_9_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_9_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_9_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_9_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_9_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_9_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_9_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_9_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_9_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_9_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_9_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_9_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_9_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_9_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_9_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_9_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_9_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_9_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_9_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_9_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_9_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_9_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_9_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_9_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_9_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_9_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_9_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_9_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_9_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_9_io_to_pes_14_in_bits),
    .io_to_mem_valid(PENetwork_9_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_9_io_to_mem_bits)
  );
  PENetwork PENetwork_10 ( // @[pe.scala 227:13]
    .io_to_pes_0_in_valid(PENetwork_10_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_10_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_10_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_10_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_10_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_10_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_10_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_10_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_10_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_10_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_10_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_10_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_10_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_10_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_10_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_10_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_10_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_10_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_10_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_10_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_10_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_10_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_10_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_10_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_10_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_10_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_10_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_10_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_10_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_10_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_10_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_10_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_10_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_10_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_10_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_10_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_10_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_10_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_10_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_10_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_10_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_10_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_10_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_10_io_to_pes_10_out_bits),
    .io_to_pes_11_in_valid(PENetwork_10_io_to_pes_11_in_valid),
    .io_to_pes_11_in_bits(PENetwork_10_io_to_pes_11_in_bits),
    .io_to_pes_11_out_valid(PENetwork_10_io_to_pes_11_out_valid),
    .io_to_pes_11_out_bits(PENetwork_10_io_to_pes_11_out_bits),
    .io_to_pes_12_in_valid(PENetwork_10_io_to_pes_12_in_valid),
    .io_to_pes_12_in_bits(PENetwork_10_io_to_pes_12_in_bits),
    .io_to_pes_12_out_valid(PENetwork_10_io_to_pes_12_out_valid),
    .io_to_pes_12_out_bits(PENetwork_10_io_to_pes_12_out_bits),
    .io_to_pes_13_in_valid(PENetwork_10_io_to_pes_13_in_valid),
    .io_to_pes_13_in_bits(PENetwork_10_io_to_pes_13_in_bits),
    .io_to_pes_13_out_valid(PENetwork_10_io_to_pes_13_out_valid),
    .io_to_pes_13_out_bits(PENetwork_10_io_to_pes_13_out_bits),
    .io_to_pes_14_in_valid(PENetwork_10_io_to_pes_14_in_valid),
    .io_to_pes_14_in_bits(PENetwork_10_io_to_pes_14_in_bits),
    .io_to_mem_valid(PENetwork_10_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_10_io_to_mem_bits)
  );
  PENetwork_11 PENetwork_11 ( // @[pe.scala 227:13]
    .io_to_pes_0_in_valid(PENetwork_11_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_11_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_11_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_11_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_11_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_11_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_11_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_11_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_11_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_11_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_11_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_11_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_11_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_11_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_11_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_11_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_11_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_11_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_11_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_11_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_11_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_11_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_11_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_11_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_11_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_11_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_11_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_11_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_11_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_11_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_11_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_11_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_11_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_11_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_11_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_11_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_11_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_11_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_11_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_11_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_11_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_11_io_to_pes_10_in_bits),
    .io_to_mem_valid(PENetwork_11_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_11_io_to_mem_bits)
  );
  PENetwork_11 PENetwork_12 ( // @[pe.scala 227:13]
    .io_to_pes_0_in_valid(PENetwork_12_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_12_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_12_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_12_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_12_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_12_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_12_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_12_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_12_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_12_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_12_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_12_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_12_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_12_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_12_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_12_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_12_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_12_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_12_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_12_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_12_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_12_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_12_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_12_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_12_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_12_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_12_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_12_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_12_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_12_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_12_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_12_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_12_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_12_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_12_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_12_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_12_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_12_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_12_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_12_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_12_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_12_io_to_pes_10_in_bits),
    .io_to_mem_valid(PENetwork_12_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_12_io_to_mem_bits)
  );
  PENetwork_11 PENetwork_13 ( // @[pe.scala 227:13]
    .io_to_pes_0_in_valid(PENetwork_13_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_13_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_13_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_13_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_13_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_13_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_13_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_13_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_13_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_13_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_13_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_13_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_13_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_13_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_13_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_13_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_13_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_13_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_13_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_13_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_13_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_13_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_13_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_13_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_13_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_13_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_13_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_13_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_13_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_13_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_13_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_13_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_13_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_13_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_13_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_13_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_13_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_13_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_13_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_13_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_13_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_13_io_to_pes_10_in_bits),
    .io_to_mem_valid(PENetwork_13_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_13_io_to_mem_bits)
  );
  PENetwork_11 PENetwork_14 ( // @[pe.scala 227:13]
    .io_to_pes_0_in_valid(PENetwork_14_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_14_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_14_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_14_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_14_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_14_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_14_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_14_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_14_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_14_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_14_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_14_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_14_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_14_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_14_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_14_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_14_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_14_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_14_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_14_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_14_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_14_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_14_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_14_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_14_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_14_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_14_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_14_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_14_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_14_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_14_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_14_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_14_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_14_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_14_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_14_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_14_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_14_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_14_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_14_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_14_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_14_io_to_pes_10_in_bits),
    .io_to_mem_valid(PENetwork_14_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_14_io_to_mem_bits)
  );
  PENetwork_11 PENetwork_15 ( // @[pe.scala 227:13]
    .io_to_pes_0_in_valid(PENetwork_15_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_15_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_15_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_15_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_15_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_15_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_15_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_15_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_15_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_15_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_15_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_15_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_15_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_15_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_15_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_15_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_15_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_15_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_15_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_15_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_15_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_15_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_15_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_15_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_15_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_15_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_15_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_15_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_15_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_15_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_15_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_15_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_15_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_15_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_15_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_15_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_15_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_15_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_15_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_15_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_15_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_15_io_to_pes_10_in_bits),
    .io_to_mem_valid(PENetwork_15_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_15_io_to_mem_bits)
  );
  PENetwork_11 PENetwork_16 ( // @[pe.scala 227:13]
    .io_to_pes_0_in_valid(PENetwork_16_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_16_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_16_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_16_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_16_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_16_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_16_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_16_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_16_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_16_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_16_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_16_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_16_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_16_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_16_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_16_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_16_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_16_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_16_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_16_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_16_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_16_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_16_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_16_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_16_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_16_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_16_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_16_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_16_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_16_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_16_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_16_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_16_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_16_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_16_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_16_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_16_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_16_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_16_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_16_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_16_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_16_io_to_pes_10_in_bits),
    .io_to_mem_valid(PENetwork_16_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_16_io_to_mem_bits)
  );
  PENetwork_11 PENetwork_17 ( // @[pe.scala 227:13]
    .io_to_pes_0_in_valid(PENetwork_17_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_17_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_17_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_17_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_17_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_17_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_17_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_17_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_17_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_17_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_17_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_17_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_17_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_17_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_17_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_17_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_17_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_17_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_17_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_17_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_17_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_17_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_17_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_17_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_17_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_17_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_17_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_17_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_17_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_17_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_17_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_17_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_17_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_17_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_17_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_17_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_17_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_17_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_17_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_17_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_17_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_17_io_to_pes_10_in_bits),
    .io_to_mem_valid(PENetwork_17_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_17_io_to_mem_bits)
  );
  PENetwork_11 PENetwork_18 ( // @[pe.scala 227:13]
    .io_to_pes_0_in_valid(PENetwork_18_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_18_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_18_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_18_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_18_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_18_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_18_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_18_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_18_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_18_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_18_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_18_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_18_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_18_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_18_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_18_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_18_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_18_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_18_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_18_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_18_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_18_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_18_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_18_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_18_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_18_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_18_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_18_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_18_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_18_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_18_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_18_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_18_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_18_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_18_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_18_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_18_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_18_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_18_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_18_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_18_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_18_io_to_pes_10_in_bits),
    .io_to_mem_valid(PENetwork_18_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_18_io_to_mem_bits)
  );
  PENetwork_11 PENetwork_19 ( // @[pe.scala 227:13]
    .io_to_pes_0_in_valid(PENetwork_19_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_19_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_19_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_19_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_19_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_19_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_19_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_19_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_19_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_19_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_19_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_19_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_19_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_19_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_19_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_19_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_19_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_19_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_19_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_19_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_19_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_19_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_19_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_19_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_19_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_19_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_19_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_19_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_19_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_19_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_19_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_19_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_19_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_19_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_19_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_19_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_19_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_19_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_19_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_19_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_19_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_19_io_to_pes_10_in_bits),
    .io_to_mem_valid(PENetwork_19_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_19_io_to_mem_bits)
  );
  PENetwork_11 PENetwork_20 ( // @[pe.scala 227:13]
    .io_to_pes_0_in_valid(PENetwork_20_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_20_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_20_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_20_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_20_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_20_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_20_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_20_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_20_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_20_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_20_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_20_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_20_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_20_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_20_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_20_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_20_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_20_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_20_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_20_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_20_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_20_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_20_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_20_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_20_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_20_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_20_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_20_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_20_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_20_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_20_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_20_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_20_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_20_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_20_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_20_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_20_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_20_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_20_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_20_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_20_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_20_io_to_pes_10_in_bits),
    .io_to_mem_valid(PENetwork_20_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_20_io_to_mem_bits)
  );
  PENetwork_11 PENetwork_21 ( // @[pe.scala 227:13]
    .io_to_pes_0_in_valid(PENetwork_21_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_21_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_21_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_21_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_21_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_21_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_21_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_21_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_21_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_21_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_21_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_21_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_21_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_21_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_21_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_21_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_21_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_21_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_21_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_21_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_21_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_21_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_21_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_21_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_21_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_21_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_21_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_21_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_21_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_21_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_21_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_21_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_21_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_21_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_21_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_21_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_21_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_21_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_21_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_21_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_21_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_21_io_to_pes_10_in_bits),
    .io_to_mem_valid(PENetwork_21_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_21_io_to_mem_bits)
  );
  PENetwork_11 PENetwork_22 ( // @[pe.scala 227:13]
    .io_to_pes_0_in_valid(PENetwork_22_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_22_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_22_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_22_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_22_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_22_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_22_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_22_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_22_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_22_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_22_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_22_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_22_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_22_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_22_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_22_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_22_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_22_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_22_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_22_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_22_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_22_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_22_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_22_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_22_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_22_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_22_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_22_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_22_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_22_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_22_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_22_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_22_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_22_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_22_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_22_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_22_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_22_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_22_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_22_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_22_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_22_io_to_pes_10_in_bits),
    .io_to_mem_valid(PENetwork_22_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_22_io_to_mem_bits)
  );
  PENetwork_11 PENetwork_23 ( // @[pe.scala 227:13]
    .io_to_pes_0_in_valid(PENetwork_23_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_23_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_23_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_23_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_23_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_23_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_23_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_23_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_23_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_23_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_23_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_23_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_23_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_23_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_23_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_23_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_23_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_23_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_23_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_23_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_23_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_23_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_23_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_23_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_23_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_23_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_23_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_23_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_23_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_23_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_23_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_23_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_23_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_23_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_23_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_23_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_23_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_23_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_23_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_23_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_23_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_23_io_to_pes_10_in_bits),
    .io_to_mem_valid(PENetwork_23_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_23_io_to_mem_bits)
  );
  PENetwork_11 PENetwork_24 ( // @[pe.scala 227:13]
    .io_to_pes_0_in_valid(PENetwork_24_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_24_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_24_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_24_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_24_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_24_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_24_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_24_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_24_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_24_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_24_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_24_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_24_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_24_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_24_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_24_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_24_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_24_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_24_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_24_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_24_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_24_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_24_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_24_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_24_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_24_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_24_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_24_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_24_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_24_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_24_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_24_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_24_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_24_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_24_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_24_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_24_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_24_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_24_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_24_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_24_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_24_io_to_pes_10_in_bits),
    .io_to_mem_valid(PENetwork_24_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_24_io_to_mem_bits)
  );
  PENetwork_11 PENetwork_25 ( // @[pe.scala 227:13]
    .io_to_pes_0_in_valid(PENetwork_25_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_25_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_25_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_25_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_25_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_25_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_25_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_25_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_25_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_25_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_25_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_25_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_25_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_25_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_25_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_25_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_25_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_25_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_25_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_25_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_25_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_25_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_25_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_25_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_25_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_25_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_25_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_25_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_25_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_25_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_25_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_25_io_to_pes_7_out_bits),
    .io_to_pes_8_in_valid(PENetwork_25_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_25_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_25_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_25_io_to_pes_8_out_bits),
    .io_to_pes_9_in_valid(PENetwork_25_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_25_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_25_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_25_io_to_pes_9_out_bits),
    .io_to_pes_10_in_valid(PENetwork_25_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_25_io_to_pes_10_in_bits),
    .io_to_mem_valid(PENetwork_25_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_25_io_to_mem_bits)
  );
  PENetwork_26 PENetwork_26 ( // @[pe.scala 227:13]
    .clock(PENetwork_26_clock),
    .io_to_pes_0_out_valid(PENetwork_26_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_26_io_to_pes_0_out_bits),
    .io_to_pes_0_sig_stat2trans(PENetwork_26_io_to_pes_0_sig_stat2trans),
    .io_to_pes_0_out_ready(PENetwork_26_io_to_pes_0_out_ready),
    .io_to_pes_1_in_valid(PENetwork_26_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_26_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_26_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_26_io_to_pes_1_out_bits),
    .io_to_pes_1_sig_stat2trans(PENetwork_26_io_to_pes_1_sig_stat2trans),
    .io_to_pes_1_in_ready(PENetwork_26_io_to_pes_1_in_ready),
    .io_to_pes_1_out_ready(PENetwork_26_io_to_pes_1_out_ready),
    .io_to_pes_2_in_valid(PENetwork_26_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_26_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_26_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_26_io_to_pes_2_out_bits),
    .io_to_pes_2_sig_stat2trans(PENetwork_26_io_to_pes_2_sig_stat2trans),
    .io_to_pes_2_in_ready(PENetwork_26_io_to_pes_2_in_ready),
    .io_to_pes_2_out_ready(PENetwork_26_io_to_pes_2_out_ready),
    .io_to_pes_3_in_valid(PENetwork_26_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_26_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_26_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_26_io_to_pes_3_out_bits),
    .io_to_pes_3_sig_stat2trans(PENetwork_26_io_to_pes_3_sig_stat2trans),
    .io_to_pes_3_in_ready(PENetwork_26_io_to_pes_3_in_ready),
    .io_to_pes_3_out_ready(PENetwork_26_io_to_pes_3_out_ready),
    .io_to_pes_4_in_valid(PENetwork_26_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_26_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_26_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_26_io_to_pes_4_out_bits),
    .io_to_pes_4_sig_stat2trans(PENetwork_26_io_to_pes_4_sig_stat2trans),
    .io_to_pes_4_in_ready(PENetwork_26_io_to_pes_4_in_ready),
    .io_to_pes_4_out_ready(PENetwork_26_io_to_pes_4_out_ready),
    .io_to_pes_5_in_valid(PENetwork_26_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_26_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_26_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_26_io_to_pes_5_out_bits),
    .io_to_pes_5_sig_stat2trans(PENetwork_26_io_to_pes_5_sig_stat2trans),
    .io_to_pes_5_in_ready(PENetwork_26_io_to_pes_5_in_ready),
    .io_to_pes_5_out_ready(PENetwork_26_io_to_pes_5_out_ready),
    .io_to_pes_6_in_valid(PENetwork_26_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_26_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_26_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_26_io_to_pes_6_out_bits),
    .io_to_pes_6_sig_stat2trans(PENetwork_26_io_to_pes_6_sig_stat2trans),
    .io_to_pes_6_in_ready(PENetwork_26_io_to_pes_6_in_ready),
    .io_to_pes_6_out_ready(PENetwork_26_io_to_pes_6_out_ready),
    .io_to_pes_7_in_valid(PENetwork_26_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_26_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_26_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_26_io_to_pes_7_out_bits),
    .io_to_pes_7_sig_stat2trans(PENetwork_26_io_to_pes_7_sig_stat2trans),
    .io_to_pes_7_in_ready(PENetwork_26_io_to_pes_7_in_ready),
    .io_to_pes_7_out_ready(PENetwork_26_io_to_pes_7_out_ready),
    .io_to_pes_8_in_valid(PENetwork_26_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_26_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_26_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_26_io_to_pes_8_out_bits),
    .io_to_pes_8_sig_stat2trans(PENetwork_26_io_to_pes_8_sig_stat2trans),
    .io_to_pes_8_in_ready(PENetwork_26_io_to_pes_8_in_ready),
    .io_to_pes_8_out_ready(PENetwork_26_io_to_pes_8_out_ready),
    .io_to_pes_9_in_valid(PENetwork_26_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_26_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_26_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_26_io_to_pes_9_out_bits),
    .io_to_pes_9_sig_stat2trans(PENetwork_26_io_to_pes_9_sig_stat2trans),
    .io_to_pes_9_in_ready(PENetwork_26_io_to_pes_9_in_ready),
    .io_to_pes_9_out_ready(PENetwork_26_io_to_pes_9_out_ready),
    .io_to_pes_10_in_valid(PENetwork_26_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_26_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_26_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_26_io_to_pes_10_out_bits),
    .io_to_pes_10_sig_stat2trans(PENetwork_26_io_to_pes_10_sig_stat2trans),
    .io_to_pes_10_in_ready(PENetwork_26_io_to_pes_10_in_ready),
    .io_to_mem_valid(PENetwork_26_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_26_io_to_mem_bits),
    .io_sig_stat2trans(PENetwork_26_io_sig_stat2trans)
  );
  PENetwork_26 PENetwork_27 ( // @[pe.scala 227:13]
    .clock(PENetwork_27_clock),
    .io_to_pes_0_out_valid(PENetwork_27_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_27_io_to_pes_0_out_bits),
    .io_to_pes_0_sig_stat2trans(PENetwork_27_io_to_pes_0_sig_stat2trans),
    .io_to_pes_0_out_ready(PENetwork_27_io_to_pes_0_out_ready),
    .io_to_pes_1_in_valid(PENetwork_27_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_27_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_27_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_27_io_to_pes_1_out_bits),
    .io_to_pes_1_sig_stat2trans(PENetwork_27_io_to_pes_1_sig_stat2trans),
    .io_to_pes_1_in_ready(PENetwork_27_io_to_pes_1_in_ready),
    .io_to_pes_1_out_ready(PENetwork_27_io_to_pes_1_out_ready),
    .io_to_pes_2_in_valid(PENetwork_27_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_27_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_27_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_27_io_to_pes_2_out_bits),
    .io_to_pes_2_sig_stat2trans(PENetwork_27_io_to_pes_2_sig_stat2trans),
    .io_to_pes_2_in_ready(PENetwork_27_io_to_pes_2_in_ready),
    .io_to_pes_2_out_ready(PENetwork_27_io_to_pes_2_out_ready),
    .io_to_pes_3_in_valid(PENetwork_27_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_27_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_27_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_27_io_to_pes_3_out_bits),
    .io_to_pes_3_sig_stat2trans(PENetwork_27_io_to_pes_3_sig_stat2trans),
    .io_to_pes_3_in_ready(PENetwork_27_io_to_pes_3_in_ready),
    .io_to_pes_3_out_ready(PENetwork_27_io_to_pes_3_out_ready),
    .io_to_pes_4_in_valid(PENetwork_27_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_27_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_27_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_27_io_to_pes_4_out_bits),
    .io_to_pes_4_sig_stat2trans(PENetwork_27_io_to_pes_4_sig_stat2trans),
    .io_to_pes_4_in_ready(PENetwork_27_io_to_pes_4_in_ready),
    .io_to_pes_4_out_ready(PENetwork_27_io_to_pes_4_out_ready),
    .io_to_pes_5_in_valid(PENetwork_27_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_27_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_27_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_27_io_to_pes_5_out_bits),
    .io_to_pes_5_sig_stat2trans(PENetwork_27_io_to_pes_5_sig_stat2trans),
    .io_to_pes_5_in_ready(PENetwork_27_io_to_pes_5_in_ready),
    .io_to_pes_5_out_ready(PENetwork_27_io_to_pes_5_out_ready),
    .io_to_pes_6_in_valid(PENetwork_27_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_27_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_27_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_27_io_to_pes_6_out_bits),
    .io_to_pes_6_sig_stat2trans(PENetwork_27_io_to_pes_6_sig_stat2trans),
    .io_to_pes_6_in_ready(PENetwork_27_io_to_pes_6_in_ready),
    .io_to_pes_6_out_ready(PENetwork_27_io_to_pes_6_out_ready),
    .io_to_pes_7_in_valid(PENetwork_27_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_27_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_27_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_27_io_to_pes_7_out_bits),
    .io_to_pes_7_sig_stat2trans(PENetwork_27_io_to_pes_7_sig_stat2trans),
    .io_to_pes_7_in_ready(PENetwork_27_io_to_pes_7_in_ready),
    .io_to_pes_7_out_ready(PENetwork_27_io_to_pes_7_out_ready),
    .io_to_pes_8_in_valid(PENetwork_27_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_27_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_27_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_27_io_to_pes_8_out_bits),
    .io_to_pes_8_sig_stat2trans(PENetwork_27_io_to_pes_8_sig_stat2trans),
    .io_to_pes_8_in_ready(PENetwork_27_io_to_pes_8_in_ready),
    .io_to_pes_8_out_ready(PENetwork_27_io_to_pes_8_out_ready),
    .io_to_pes_9_in_valid(PENetwork_27_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_27_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_27_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_27_io_to_pes_9_out_bits),
    .io_to_pes_9_sig_stat2trans(PENetwork_27_io_to_pes_9_sig_stat2trans),
    .io_to_pes_9_in_ready(PENetwork_27_io_to_pes_9_in_ready),
    .io_to_pes_9_out_ready(PENetwork_27_io_to_pes_9_out_ready),
    .io_to_pes_10_in_valid(PENetwork_27_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_27_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_27_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_27_io_to_pes_10_out_bits),
    .io_to_pes_10_sig_stat2trans(PENetwork_27_io_to_pes_10_sig_stat2trans),
    .io_to_pes_10_in_ready(PENetwork_27_io_to_pes_10_in_ready),
    .io_to_mem_valid(PENetwork_27_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_27_io_to_mem_bits),
    .io_sig_stat2trans(PENetwork_27_io_sig_stat2trans)
  );
  PENetwork_26 PENetwork_28 ( // @[pe.scala 227:13]
    .clock(PENetwork_28_clock),
    .io_to_pes_0_out_valid(PENetwork_28_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_28_io_to_pes_0_out_bits),
    .io_to_pes_0_sig_stat2trans(PENetwork_28_io_to_pes_0_sig_stat2trans),
    .io_to_pes_0_out_ready(PENetwork_28_io_to_pes_0_out_ready),
    .io_to_pes_1_in_valid(PENetwork_28_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_28_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_28_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_28_io_to_pes_1_out_bits),
    .io_to_pes_1_sig_stat2trans(PENetwork_28_io_to_pes_1_sig_stat2trans),
    .io_to_pes_1_in_ready(PENetwork_28_io_to_pes_1_in_ready),
    .io_to_pes_1_out_ready(PENetwork_28_io_to_pes_1_out_ready),
    .io_to_pes_2_in_valid(PENetwork_28_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_28_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_28_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_28_io_to_pes_2_out_bits),
    .io_to_pes_2_sig_stat2trans(PENetwork_28_io_to_pes_2_sig_stat2trans),
    .io_to_pes_2_in_ready(PENetwork_28_io_to_pes_2_in_ready),
    .io_to_pes_2_out_ready(PENetwork_28_io_to_pes_2_out_ready),
    .io_to_pes_3_in_valid(PENetwork_28_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_28_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_28_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_28_io_to_pes_3_out_bits),
    .io_to_pes_3_sig_stat2trans(PENetwork_28_io_to_pes_3_sig_stat2trans),
    .io_to_pes_3_in_ready(PENetwork_28_io_to_pes_3_in_ready),
    .io_to_pes_3_out_ready(PENetwork_28_io_to_pes_3_out_ready),
    .io_to_pes_4_in_valid(PENetwork_28_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_28_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_28_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_28_io_to_pes_4_out_bits),
    .io_to_pes_4_sig_stat2trans(PENetwork_28_io_to_pes_4_sig_stat2trans),
    .io_to_pes_4_in_ready(PENetwork_28_io_to_pes_4_in_ready),
    .io_to_pes_4_out_ready(PENetwork_28_io_to_pes_4_out_ready),
    .io_to_pes_5_in_valid(PENetwork_28_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_28_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_28_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_28_io_to_pes_5_out_bits),
    .io_to_pes_5_sig_stat2trans(PENetwork_28_io_to_pes_5_sig_stat2trans),
    .io_to_pes_5_in_ready(PENetwork_28_io_to_pes_5_in_ready),
    .io_to_pes_5_out_ready(PENetwork_28_io_to_pes_5_out_ready),
    .io_to_pes_6_in_valid(PENetwork_28_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_28_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_28_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_28_io_to_pes_6_out_bits),
    .io_to_pes_6_sig_stat2trans(PENetwork_28_io_to_pes_6_sig_stat2trans),
    .io_to_pes_6_in_ready(PENetwork_28_io_to_pes_6_in_ready),
    .io_to_pes_6_out_ready(PENetwork_28_io_to_pes_6_out_ready),
    .io_to_pes_7_in_valid(PENetwork_28_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_28_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_28_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_28_io_to_pes_7_out_bits),
    .io_to_pes_7_sig_stat2trans(PENetwork_28_io_to_pes_7_sig_stat2trans),
    .io_to_pes_7_in_ready(PENetwork_28_io_to_pes_7_in_ready),
    .io_to_pes_7_out_ready(PENetwork_28_io_to_pes_7_out_ready),
    .io_to_pes_8_in_valid(PENetwork_28_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_28_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_28_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_28_io_to_pes_8_out_bits),
    .io_to_pes_8_sig_stat2trans(PENetwork_28_io_to_pes_8_sig_stat2trans),
    .io_to_pes_8_in_ready(PENetwork_28_io_to_pes_8_in_ready),
    .io_to_pes_8_out_ready(PENetwork_28_io_to_pes_8_out_ready),
    .io_to_pes_9_in_valid(PENetwork_28_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_28_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_28_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_28_io_to_pes_9_out_bits),
    .io_to_pes_9_sig_stat2trans(PENetwork_28_io_to_pes_9_sig_stat2trans),
    .io_to_pes_9_in_ready(PENetwork_28_io_to_pes_9_in_ready),
    .io_to_pes_9_out_ready(PENetwork_28_io_to_pes_9_out_ready),
    .io_to_pes_10_in_valid(PENetwork_28_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_28_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_28_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_28_io_to_pes_10_out_bits),
    .io_to_pes_10_sig_stat2trans(PENetwork_28_io_to_pes_10_sig_stat2trans),
    .io_to_pes_10_in_ready(PENetwork_28_io_to_pes_10_in_ready),
    .io_to_mem_valid(PENetwork_28_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_28_io_to_mem_bits),
    .io_sig_stat2trans(PENetwork_28_io_sig_stat2trans)
  );
  PENetwork_26 PENetwork_29 ( // @[pe.scala 227:13]
    .clock(PENetwork_29_clock),
    .io_to_pes_0_out_valid(PENetwork_29_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_29_io_to_pes_0_out_bits),
    .io_to_pes_0_sig_stat2trans(PENetwork_29_io_to_pes_0_sig_stat2trans),
    .io_to_pes_0_out_ready(PENetwork_29_io_to_pes_0_out_ready),
    .io_to_pes_1_in_valid(PENetwork_29_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_29_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_29_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_29_io_to_pes_1_out_bits),
    .io_to_pes_1_sig_stat2trans(PENetwork_29_io_to_pes_1_sig_stat2trans),
    .io_to_pes_1_in_ready(PENetwork_29_io_to_pes_1_in_ready),
    .io_to_pes_1_out_ready(PENetwork_29_io_to_pes_1_out_ready),
    .io_to_pes_2_in_valid(PENetwork_29_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_29_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_29_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_29_io_to_pes_2_out_bits),
    .io_to_pes_2_sig_stat2trans(PENetwork_29_io_to_pes_2_sig_stat2trans),
    .io_to_pes_2_in_ready(PENetwork_29_io_to_pes_2_in_ready),
    .io_to_pes_2_out_ready(PENetwork_29_io_to_pes_2_out_ready),
    .io_to_pes_3_in_valid(PENetwork_29_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_29_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_29_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_29_io_to_pes_3_out_bits),
    .io_to_pes_3_sig_stat2trans(PENetwork_29_io_to_pes_3_sig_stat2trans),
    .io_to_pes_3_in_ready(PENetwork_29_io_to_pes_3_in_ready),
    .io_to_pes_3_out_ready(PENetwork_29_io_to_pes_3_out_ready),
    .io_to_pes_4_in_valid(PENetwork_29_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_29_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_29_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_29_io_to_pes_4_out_bits),
    .io_to_pes_4_sig_stat2trans(PENetwork_29_io_to_pes_4_sig_stat2trans),
    .io_to_pes_4_in_ready(PENetwork_29_io_to_pes_4_in_ready),
    .io_to_pes_4_out_ready(PENetwork_29_io_to_pes_4_out_ready),
    .io_to_pes_5_in_valid(PENetwork_29_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_29_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_29_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_29_io_to_pes_5_out_bits),
    .io_to_pes_5_sig_stat2trans(PENetwork_29_io_to_pes_5_sig_stat2trans),
    .io_to_pes_5_in_ready(PENetwork_29_io_to_pes_5_in_ready),
    .io_to_pes_5_out_ready(PENetwork_29_io_to_pes_5_out_ready),
    .io_to_pes_6_in_valid(PENetwork_29_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_29_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_29_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_29_io_to_pes_6_out_bits),
    .io_to_pes_6_sig_stat2trans(PENetwork_29_io_to_pes_6_sig_stat2trans),
    .io_to_pes_6_in_ready(PENetwork_29_io_to_pes_6_in_ready),
    .io_to_pes_6_out_ready(PENetwork_29_io_to_pes_6_out_ready),
    .io_to_pes_7_in_valid(PENetwork_29_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_29_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_29_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_29_io_to_pes_7_out_bits),
    .io_to_pes_7_sig_stat2trans(PENetwork_29_io_to_pes_7_sig_stat2trans),
    .io_to_pes_7_in_ready(PENetwork_29_io_to_pes_7_in_ready),
    .io_to_pes_7_out_ready(PENetwork_29_io_to_pes_7_out_ready),
    .io_to_pes_8_in_valid(PENetwork_29_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_29_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_29_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_29_io_to_pes_8_out_bits),
    .io_to_pes_8_sig_stat2trans(PENetwork_29_io_to_pes_8_sig_stat2trans),
    .io_to_pes_8_in_ready(PENetwork_29_io_to_pes_8_in_ready),
    .io_to_pes_8_out_ready(PENetwork_29_io_to_pes_8_out_ready),
    .io_to_pes_9_in_valid(PENetwork_29_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_29_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_29_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_29_io_to_pes_9_out_bits),
    .io_to_pes_9_sig_stat2trans(PENetwork_29_io_to_pes_9_sig_stat2trans),
    .io_to_pes_9_in_ready(PENetwork_29_io_to_pes_9_in_ready),
    .io_to_pes_9_out_ready(PENetwork_29_io_to_pes_9_out_ready),
    .io_to_pes_10_in_valid(PENetwork_29_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_29_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_29_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_29_io_to_pes_10_out_bits),
    .io_to_pes_10_sig_stat2trans(PENetwork_29_io_to_pes_10_sig_stat2trans),
    .io_to_pes_10_in_ready(PENetwork_29_io_to_pes_10_in_ready),
    .io_to_mem_valid(PENetwork_29_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_29_io_to_mem_bits),
    .io_sig_stat2trans(PENetwork_29_io_sig_stat2trans)
  );
  PENetwork_26 PENetwork_30 ( // @[pe.scala 227:13]
    .clock(PENetwork_30_clock),
    .io_to_pes_0_out_valid(PENetwork_30_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_30_io_to_pes_0_out_bits),
    .io_to_pes_0_sig_stat2trans(PENetwork_30_io_to_pes_0_sig_stat2trans),
    .io_to_pes_0_out_ready(PENetwork_30_io_to_pes_0_out_ready),
    .io_to_pes_1_in_valid(PENetwork_30_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_30_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_30_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_30_io_to_pes_1_out_bits),
    .io_to_pes_1_sig_stat2trans(PENetwork_30_io_to_pes_1_sig_stat2trans),
    .io_to_pes_1_in_ready(PENetwork_30_io_to_pes_1_in_ready),
    .io_to_pes_1_out_ready(PENetwork_30_io_to_pes_1_out_ready),
    .io_to_pes_2_in_valid(PENetwork_30_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_30_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_30_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_30_io_to_pes_2_out_bits),
    .io_to_pes_2_sig_stat2trans(PENetwork_30_io_to_pes_2_sig_stat2trans),
    .io_to_pes_2_in_ready(PENetwork_30_io_to_pes_2_in_ready),
    .io_to_pes_2_out_ready(PENetwork_30_io_to_pes_2_out_ready),
    .io_to_pes_3_in_valid(PENetwork_30_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_30_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_30_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_30_io_to_pes_3_out_bits),
    .io_to_pes_3_sig_stat2trans(PENetwork_30_io_to_pes_3_sig_stat2trans),
    .io_to_pes_3_in_ready(PENetwork_30_io_to_pes_3_in_ready),
    .io_to_pes_3_out_ready(PENetwork_30_io_to_pes_3_out_ready),
    .io_to_pes_4_in_valid(PENetwork_30_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_30_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_30_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_30_io_to_pes_4_out_bits),
    .io_to_pes_4_sig_stat2trans(PENetwork_30_io_to_pes_4_sig_stat2trans),
    .io_to_pes_4_in_ready(PENetwork_30_io_to_pes_4_in_ready),
    .io_to_pes_4_out_ready(PENetwork_30_io_to_pes_4_out_ready),
    .io_to_pes_5_in_valid(PENetwork_30_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_30_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_30_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_30_io_to_pes_5_out_bits),
    .io_to_pes_5_sig_stat2trans(PENetwork_30_io_to_pes_5_sig_stat2trans),
    .io_to_pes_5_in_ready(PENetwork_30_io_to_pes_5_in_ready),
    .io_to_pes_5_out_ready(PENetwork_30_io_to_pes_5_out_ready),
    .io_to_pes_6_in_valid(PENetwork_30_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_30_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_30_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_30_io_to_pes_6_out_bits),
    .io_to_pes_6_sig_stat2trans(PENetwork_30_io_to_pes_6_sig_stat2trans),
    .io_to_pes_6_in_ready(PENetwork_30_io_to_pes_6_in_ready),
    .io_to_pes_6_out_ready(PENetwork_30_io_to_pes_6_out_ready),
    .io_to_pes_7_in_valid(PENetwork_30_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_30_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_30_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_30_io_to_pes_7_out_bits),
    .io_to_pes_7_sig_stat2trans(PENetwork_30_io_to_pes_7_sig_stat2trans),
    .io_to_pes_7_in_ready(PENetwork_30_io_to_pes_7_in_ready),
    .io_to_pes_7_out_ready(PENetwork_30_io_to_pes_7_out_ready),
    .io_to_pes_8_in_valid(PENetwork_30_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_30_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_30_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_30_io_to_pes_8_out_bits),
    .io_to_pes_8_sig_stat2trans(PENetwork_30_io_to_pes_8_sig_stat2trans),
    .io_to_pes_8_in_ready(PENetwork_30_io_to_pes_8_in_ready),
    .io_to_pes_8_out_ready(PENetwork_30_io_to_pes_8_out_ready),
    .io_to_pes_9_in_valid(PENetwork_30_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_30_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_30_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_30_io_to_pes_9_out_bits),
    .io_to_pes_9_sig_stat2trans(PENetwork_30_io_to_pes_9_sig_stat2trans),
    .io_to_pes_9_in_ready(PENetwork_30_io_to_pes_9_in_ready),
    .io_to_pes_9_out_ready(PENetwork_30_io_to_pes_9_out_ready),
    .io_to_pes_10_in_valid(PENetwork_30_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_30_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_30_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_30_io_to_pes_10_out_bits),
    .io_to_pes_10_sig_stat2trans(PENetwork_30_io_to_pes_10_sig_stat2trans),
    .io_to_pes_10_in_ready(PENetwork_30_io_to_pes_10_in_ready),
    .io_to_mem_valid(PENetwork_30_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_30_io_to_mem_bits),
    .io_sig_stat2trans(PENetwork_30_io_sig_stat2trans)
  );
  PENetwork_26 PENetwork_31 ( // @[pe.scala 227:13]
    .clock(PENetwork_31_clock),
    .io_to_pes_0_out_valid(PENetwork_31_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_31_io_to_pes_0_out_bits),
    .io_to_pes_0_sig_stat2trans(PENetwork_31_io_to_pes_0_sig_stat2trans),
    .io_to_pes_0_out_ready(PENetwork_31_io_to_pes_0_out_ready),
    .io_to_pes_1_in_valid(PENetwork_31_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_31_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_31_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_31_io_to_pes_1_out_bits),
    .io_to_pes_1_sig_stat2trans(PENetwork_31_io_to_pes_1_sig_stat2trans),
    .io_to_pes_1_in_ready(PENetwork_31_io_to_pes_1_in_ready),
    .io_to_pes_1_out_ready(PENetwork_31_io_to_pes_1_out_ready),
    .io_to_pes_2_in_valid(PENetwork_31_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_31_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_31_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_31_io_to_pes_2_out_bits),
    .io_to_pes_2_sig_stat2trans(PENetwork_31_io_to_pes_2_sig_stat2trans),
    .io_to_pes_2_in_ready(PENetwork_31_io_to_pes_2_in_ready),
    .io_to_pes_2_out_ready(PENetwork_31_io_to_pes_2_out_ready),
    .io_to_pes_3_in_valid(PENetwork_31_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_31_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_31_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_31_io_to_pes_3_out_bits),
    .io_to_pes_3_sig_stat2trans(PENetwork_31_io_to_pes_3_sig_stat2trans),
    .io_to_pes_3_in_ready(PENetwork_31_io_to_pes_3_in_ready),
    .io_to_pes_3_out_ready(PENetwork_31_io_to_pes_3_out_ready),
    .io_to_pes_4_in_valid(PENetwork_31_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_31_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_31_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_31_io_to_pes_4_out_bits),
    .io_to_pes_4_sig_stat2trans(PENetwork_31_io_to_pes_4_sig_stat2trans),
    .io_to_pes_4_in_ready(PENetwork_31_io_to_pes_4_in_ready),
    .io_to_pes_4_out_ready(PENetwork_31_io_to_pes_4_out_ready),
    .io_to_pes_5_in_valid(PENetwork_31_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_31_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_31_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_31_io_to_pes_5_out_bits),
    .io_to_pes_5_sig_stat2trans(PENetwork_31_io_to_pes_5_sig_stat2trans),
    .io_to_pes_5_in_ready(PENetwork_31_io_to_pes_5_in_ready),
    .io_to_pes_5_out_ready(PENetwork_31_io_to_pes_5_out_ready),
    .io_to_pes_6_in_valid(PENetwork_31_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_31_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_31_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_31_io_to_pes_6_out_bits),
    .io_to_pes_6_sig_stat2trans(PENetwork_31_io_to_pes_6_sig_stat2trans),
    .io_to_pes_6_in_ready(PENetwork_31_io_to_pes_6_in_ready),
    .io_to_pes_6_out_ready(PENetwork_31_io_to_pes_6_out_ready),
    .io_to_pes_7_in_valid(PENetwork_31_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_31_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_31_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_31_io_to_pes_7_out_bits),
    .io_to_pes_7_sig_stat2trans(PENetwork_31_io_to_pes_7_sig_stat2trans),
    .io_to_pes_7_in_ready(PENetwork_31_io_to_pes_7_in_ready),
    .io_to_pes_7_out_ready(PENetwork_31_io_to_pes_7_out_ready),
    .io_to_pes_8_in_valid(PENetwork_31_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_31_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_31_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_31_io_to_pes_8_out_bits),
    .io_to_pes_8_sig_stat2trans(PENetwork_31_io_to_pes_8_sig_stat2trans),
    .io_to_pes_8_in_ready(PENetwork_31_io_to_pes_8_in_ready),
    .io_to_pes_8_out_ready(PENetwork_31_io_to_pes_8_out_ready),
    .io_to_pes_9_in_valid(PENetwork_31_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_31_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_31_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_31_io_to_pes_9_out_bits),
    .io_to_pes_9_sig_stat2trans(PENetwork_31_io_to_pes_9_sig_stat2trans),
    .io_to_pes_9_in_ready(PENetwork_31_io_to_pes_9_in_ready),
    .io_to_pes_9_out_ready(PENetwork_31_io_to_pes_9_out_ready),
    .io_to_pes_10_in_valid(PENetwork_31_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_31_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_31_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_31_io_to_pes_10_out_bits),
    .io_to_pes_10_sig_stat2trans(PENetwork_31_io_to_pes_10_sig_stat2trans),
    .io_to_pes_10_in_ready(PENetwork_31_io_to_pes_10_in_ready),
    .io_to_mem_valid(PENetwork_31_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_31_io_to_mem_bits),
    .io_sig_stat2trans(PENetwork_31_io_sig_stat2trans)
  );
  PENetwork_26 PENetwork_32 ( // @[pe.scala 227:13]
    .clock(PENetwork_32_clock),
    .io_to_pes_0_out_valid(PENetwork_32_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_32_io_to_pes_0_out_bits),
    .io_to_pes_0_sig_stat2trans(PENetwork_32_io_to_pes_0_sig_stat2trans),
    .io_to_pes_0_out_ready(PENetwork_32_io_to_pes_0_out_ready),
    .io_to_pes_1_in_valid(PENetwork_32_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_32_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_32_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_32_io_to_pes_1_out_bits),
    .io_to_pes_1_sig_stat2trans(PENetwork_32_io_to_pes_1_sig_stat2trans),
    .io_to_pes_1_in_ready(PENetwork_32_io_to_pes_1_in_ready),
    .io_to_pes_1_out_ready(PENetwork_32_io_to_pes_1_out_ready),
    .io_to_pes_2_in_valid(PENetwork_32_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_32_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_32_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_32_io_to_pes_2_out_bits),
    .io_to_pes_2_sig_stat2trans(PENetwork_32_io_to_pes_2_sig_stat2trans),
    .io_to_pes_2_in_ready(PENetwork_32_io_to_pes_2_in_ready),
    .io_to_pes_2_out_ready(PENetwork_32_io_to_pes_2_out_ready),
    .io_to_pes_3_in_valid(PENetwork_32_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_32_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_32_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_32_io_to_pes_3_out_bits),
    .io_to_pes_3_sig_stat2trans(PENetwork_32_io_to_pes_3_sig_stat2trans),
    .io_to_pes_3_in_ready(PENetwork_32_io_to_pes_3_in_ready),
    .io_to_pes_3_out_ready(PENetwork_32_io_to_pes_3_out_ready),
    .io_to_pes_4_in_valid(PENetwork_32_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_32_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_32_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_32_io_to_pes_4_out_bits),
    .io_to_pes_4_sig_stat2trans(PENetwork_32_io_to_pes_4_sig_stat2trans),
    .io_to_pes_4_in_ready(PENetwork_32_io_to_pes_4_in_ready),
    .io_to_pes_4_out_ready(PENetwork_32_io_to_pes_4_out_ready),
    .io_to_pes_5_in_valid(PENetwork_32_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_32_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_32_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_32_io_to_pes_5_out_bits),
    .io_to_pes_5_sig_stat2trans(PENetwork_32_io_to_pes_5_sig_stat2trans),
    .io_to_pes_5_in_ready(PENetwork_32_io_to_pes_5_in_ready),
    .io_to_pes_5_out_ready(PENetwork_32_io_to_pes_5_out_ready),
    .io_to_pes_6_in_valid(PENetwork_32_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_32_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_32_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_32_io_to_pes_6_out_bits),
    .io_to_pes_6_sig_stat2trans(PENetwork_32_io_to_pes_6_sig_stat2trans),
    .io_to_pes_6_in_ready(PENetwork_32_io_to_pes_6_in_ready),
    .io_to_pes_6_out_ready(PENetwork_32_io_to_pes_6_out_ready),
    .io_to_pes_7_in_valid(PENetwork_32_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_32_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_32_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_32_io_to_pes_7_out_bits),
    .io_to_pes_7_sig_stat2trans(PENetwork_32_io_to_pes_7_sig_stat2trans),
    .io_to_pes_7_in_ready(PENetwork_32_io_to_pes_7_in_ready),
    .io_to_pes_7_out_ready(PENetwork_32_io_to_pes_7_out_ready),
    .io_to_pes_8_in_valid(PENetwork_32_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_32_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_32_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_32_io_to_pes_8_out_bits),
    .io_to_pes_8_sig_stat2trans(PENetwork_32_io_to_pes_8_sig_stat2trans),
    .io_to_pes_8_in_ready(PENetwork_32_io_to_pes_8_in_ready),
    .io_to_pes_8_out_ready(PENetwork_32_io_to_pes_8_out_ready),
    .io_to_pes_9_in_valid(PENetwork_32_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_32_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_32_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_32_io_to_pes_9_out_bits),
    .io_to_pes_9_sig_stat2trans(PENetwork_32_io_to_pes_9_sig_stat2trans),
    .io_to_pes_9_in_ready(PENetwork_32_io_to_pes_9_in_ready),
    .io_to_pes_9_out_ready(PENetwork_32_io_to_pes_9_out_ready),
    .io_to_pes_10_in_valid(PENetwork_32_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_32_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_32_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_32_io_to_pes_10_out_bits),
    .io_to_pes_10_sig_stat2trans(PENetwork_32_io_to_pes_10_sig_stat2trans),
    .io_to_pes_10_in_ready(PENetwork_32_io_to_pes_10_in_ready),
    .io_to_mem_valid(PENetwork_32_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_32_io_to_mem_bits),
    .io_sig_stat2trans(PENetwork_32_io_sig_stat2trans)
  );
  PENetwork_26 PENetwork_33 ( // @[pe.scala 227:13]
    .clock(PENetwork_33_clock),
    .io_to_pes_0_out_valid(PENetwork_33_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_33_io_to_pes_0_out_bits),
    .io_to_pes_0_sig_stat2trans(PENetwork_33_io_to_pes_0_sig_stat2trans),
    .io_to_pes_0_out_ready(PENetwork_33_io_to_pes_0_out_ready),
    .io_to_pes_1_in_valid(PENetwork_33_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_33_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_33_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_33_io_to_pes_1_out_bits),
    .io_to_pes_1_sig_stat2trans(PENetwork_33_io_to_pes_1_sig_stat2trans),
    .io_to_pes_1_in_ready(PENetwork_33_io_to_pes_1_in_ready),
    .io_to_pes_1_out_ready(PENetwork_33_io_to_pes_1_out_ready),
    .io_to_pes_2_in_valid(PENetwork_33_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_33_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_33_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_33_io_to_pes_2_out_bits),
    .io_to_pes_2_sig_stat2trans(PENetwork_33_io_to_pes_2_sig_stat2trans),
    .io_to_pes_2_in_ready(PENetwork_33_io_to_pes_2_in_ready),
    .io_to_pes_2_out_ready(PENetwork_33_io_to_pes_2_out_ready),
    .io_to_pes_3_in_valid(PENetwork_33_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_33_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_33_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_33_io_to_pes_3_out_bits),
    .io_to_pes_3_sig_stat2trans(PENetwork_33_io_to_pes_3_sig_stat2trans),
    .io_to_pes_3_in_ready(PENetwork_33_io_to_pes_3_in_ready),
    .io_to_pes_3_out_ready(PENetwork_33_io_to_pes_3_out_ready),
    .io_to_pes_4_in_valid(PENetwork_33_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_33_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_33_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_33_io_to_pes_4_out_bits),
    .io_to_pes_4_sig_stat2trans(PENetwork_33_io_to_pes_4_sig_stat2trans),
    .io_to_pes_4_in_ready(PENetwork_33_io_to_pes_4_in_ready),
    .io_to_pes_4_out_ready(PENetwork_33_io_to_pes_4_out_ready),
    .io_to_pes_5_in_valid(PENetwork_33_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_33_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_33_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_33_io_to_pes_5_out_bits),
    .io_to_pes_5_sig_stat2trans(PENetwork_33_io_to_pes_5_sig_stat2trans),
    .io_to_pes_5_in_ready(PENetwork_33_io_to_pes_5_in_ready),
    .io_to_pes_5_out_ready(PENetwork_33_io_to_pes_5_out_ready),
    .io_to_pes_6_in_valid(PENetwork_33_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_33_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_33_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_33_io_to_pes_6_out_bits),
    .io_to_pes_6_sig_stat2trans(PENetwork_33_io_to_pes_6_sig_stat2trans),
    .io_to_pes_6_in_ready(PENetwork_33_io_to_pes_6_in_ready),
    .io_to_pes_6_out_ready(PENetwork_33_io_to_pes_6_out_ready),
    .io_to_pes_7_in_valid(PENetwork_33_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_33_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_33_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_33_io_to_pes_7_out_bits),
    .io_to_pes_7_sig_stat2trans(PENetwork_33_io_to_pes_7_sig_stat2trans),
    .io_to_pes_7_in_ready(PENetwork_33_io_to_pes_7_in_ready),
    .io_to_pes_7_out_ready(PENetwork_33_io_to_pes_7_out_ready),
    .io_to_pes_8_in_valid(PENetwork_33_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_33_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_33_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_33_io_to_pes_8_out_bits),
    .io_to_pes_8_sig_stat2trans(PENetwork_33_io_to_pes_8_sig_stat2trans),
    .io_to_pes_8_in_ready(PENetwork_33_io_to_pes_8_in_ready),
    .io_to_pes_8_out_ready(PENetwork_33_io_to_pes_8_out_ready),
    .io_to_pes_9_in_valid(PENetwork_33_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_33_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_33_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_33_io_to_pes_9_out_bits),
    .io_to_pes_9_sig_stat2trans(PENetwork_33_io_to_pes_9_sig_stat2trans),
    .io_to_pes_9_in_ready(PENetwork_33_io_to_pes_9_in_ready),
    .io_to_pes_9_out_ready(PENetwork_33_io_to_pes_9_out_ready),
    .io_to_pes_10_in_valid(PENetwork_33_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_33_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_33_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_33_io_to_pes_10_out_bits),
    .io_to_pes_10_sig_stat2trans(PENetwork_33_io_to_pes_10_sig_stat2trans),
    .io_to_pes_10_in_ready(PENetwork_33_io_to_pes_10_in_ready),
    .io_to_mem_valid(PENetwork_33_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_33_io_to_mem_bits),
    .io_sig_stat2trans(PENetwork_33_io_sig_stat2trans)
  );
  PENetwork_26 PENetwork_34 ( // @[pe.scala 227:13]
    .clock(PENetwork_34_clock),
    .io_to_pes_0_out_valid(PENetwork_34_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_34_io_to_pes_0_out_bits),
    .io_to_pes_0_sig_stat2trans(PENetwork_34_io_to_pes_0_sig_stat2trans),
    .io_to_pes_0_out_ready(PENetwork_34_io_to_pes_0_out_ready),
    .io_to_pes_1_in_valid(PENetwork_34_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_34_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_34_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_34_io_to_pes_1_out_bits),
    .io_to_pes_1_sig_stat2trans(PENetwork_34_io_to_pes_1_sig_stat2trans),
    .io_to_pes_1_in_ready(PENetwork_34_io_to_pes_1_in_ready),
    .io_to_pes_1_out_ready(PENetwork_34_io_to_pes_1_out_ready),
    .io_to_pes_2_in_valid(PENetwork_34_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_34_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_34_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_34_io_to_pes_2_out_bits),
    .io_to_pes_2_sig_stat2trans(PENetwork_34_io_to_pes_2_sig_stat2trans),
    .io_to_pes_2_in_ready(PENetwork_34_io_to_pes_2_in_ready),
    .io_to_pes_2_out_ready(PENetwork_34_io_to_pes_2_out_ready),
    .io_to_pes_3_in_valid(PENetwork_34_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_34_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_34_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_34_io_to_pes_3_out_bits),
    .io_to_pes_3_sig_stat2trans(PENetwork_34_io_to_pes_3_sig_stat2trans),
    .io_to_pes_3_in_ready(PENetwork_34_io_to_pes_3_in_ready),
    .io_to_pes_3_out_ready(PENetwork_34_io_to_pes_3_out_ready),
    .io_to_pes_4_in_valid(PENetwork_34_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_34_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_34_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_34_io_to_pes_4_out_bits),
    .io_to_pes_4_sig_stat2trans(PENetwork_34_io_to_pes_4_sig_stat2trans),
    .io_to_pes_4_in_ready(PENetwork_34_io_to_pes_4_in_ready),
    .io_to_pes_4_out_ready(PENetwork_34_io_to_pes_4_out_ready),
    .io_to_pes_5_in_valid(PENetwork_34_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_34_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_34_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_34_io_to_pes_5_out_bits),
    .io_to_pes_5_sig_stat2trans(PENetwork_34_io_to_pes_5_sig_stat2trans),
    .io_to_pes_5_in_ready(PENetwork_34_io_to_pes_5_in_ready),
    .io_to_pes_5_out_ready(PENetwork_34_io_to_pes_5_out_ready),
    .io_to_pes_6_in_valid(PENetwork_34_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_34_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_34_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_34_io_to_pes_6_out_bits),
    .io_to_pes_6_sig_stat2trans(PENetwork_34_io_to_pes_6_sig_stat2trans),
    .io_to_pes_6_in_ready(PENetwork_34_io_to_pes_6_in_ready),
    .io_to_pes_6_out_ready(PENetwork_34_io_to_pes_6_out_ready),
    .io_to_pes_7_in_valid(PENetwork_34_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_34_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_34_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_34_io_to_pes_7_out_bits),
    .io_to_pes_7_sig_stat2trans(PENetwork_34_io_to_pes_7_sig_stat2trans),
    .io_to_pes_7_in_ready(PENetwork_34_io_to_pes_7_in_ready),
    .io_to_pes_7_out_ready(PENetwork_34_io_to_pes_7_out_ready),
    .io_to_pes_8_in_valid(PENetwork_34_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_34_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_34_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_34_io_to_pes_8_out_bits),
    .io_to_pes_8_sig_stat2trans(PENetwork_34_io_to_pes_8_sig_stat2trans),
    .io_to_pes_8_in_ready(PENetwork_34_io_to_pes_8_in_ready),
    .io_to_pes_8_out_ready(PENetwork_34_io_to_pes_8_out_ready),
    .io_to_pes_9_in_valid(PENetwork_34_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_34_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_34_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_34_io_to_pes_9_out_bits),
    .io_to_pes_9_sig_stat2trans(PENetwork_34_io_to_pes_9_sig_stat2trans),
    .io_to_pes_9_in_ready(PENetwork_34_io_to_pes_9_in_ready),
    .io_to_pes_9_out_ready(PENetwork_34_io_to_pes_9_out_ready),
    .io_to_pes_10_in_valid(PENetwork_34_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_34_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_34_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_34_io_to_pes_10_out_bits),
    .io_to_pes_10_sig_stat2trans(PENetwork_34_io_to_pes_10_sig_stat2trans),
    .io_to_pes_10_in_ready(PENetwork_34_io_to_pes_10_in_ready),
    .io_to_mem_valid(PENetwork_34_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_34_io_to_mem_bits),
    .io_sig_stat2trans(PENetwork_34_io_sig_stat2trans)
  );
  PENetwork_26 PENetwork_35 ( // @[pe.scala 227:13]
    .clock(PENetwork_35_clock),
    .io_to_pes_0_out_valid(PENetwork_35_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_35_io_to_pes_0_out_bits),
    .io_to_pes_0_sig_stat2trans(PENetwork_35_io_to_pes_0_sig_stat2trans),
    .io_to_pes_0_out_ready(PENetwork_35_io_to_pes_0_out_ready),
    .io_to_pes_1_in_valid(PENetwork_35_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_35_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_35_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_35_io_to_pes_1_out_bits),
    .io_to_pes_1_sig_stat2trans(PENetwork_35_io_to_pes_1_sig_stat2trans),
    .io_to_pes_1_in_ready(PENetwork_35_io_to_pes_1_in_ready),
    .io_to_pes_1_out_ready(PENetwork_35_io_to_pes_1_out_ready),
    .io_to_pes_2_in_valid(PENetwork_35_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_35_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_35_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_35_io_to_pes_2_out_bits),
    .io_to_pes_2_sig_stat2trans(PENetwork_35_io_to_pes_2_sig_stat2trans),
    .io_to_pes_2_in_ready(PENetwork_35_io_to_pes_2_in_ready),
    .io_to_pes_2_out_ready(PENetwork_35_io_to_pes_2_out_ready),
    .io_to_pes_3_in_valid(PENetwork_35_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_35_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_35_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_35_io_to_pes_3_out_bits),
    .io_to_pes_3_sig_stat2trans(PENetwork_35_io_to_pes_3_sig_stat2trans),
    .io_to_pes_3_in_ready(PENetwork_35_io_to_pes_3_in_ready),
    .io_to_pes_3_out_ready(PENetwork_35_io_to_pes_3_out_ready),
    .io_to_pes_4_in_valid(PENetwork_35_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_35_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_35_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_35_io_to_pes_4_out_bits),
    .io_to_pes_4_sig_stat2trans(PENetwork_35_io_to_pes_4_sig_stat2trans),
    .io_to_pes_4_in_ready(PENetwork_35_io_to_pes_4_in_ready),
    .io_to_pes_4_out_ready(PENetwork_35_io_to_pes_4_out_ready),
    .io_to_pes_5_in_valid(PENetwork_35_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_35_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_35_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_35_io_to_pes_5_out_bits),
    .io_to_pes_5_sig_stat2trans(PENetwork_35_io_to_pes_5_sig_stat2trans),
    .io_to_pes_5_in_ready(PENetwork_35_io_to_pes_5_in_ready),
    .io_to_pes_5_out_ready(PENetwork_35_io_to_pes_5_out_ready),
    .io_to_pes_6_in_valid(PENetwork_35_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_35_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_35_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_35_io_to_pes_6_out_bits),
    .io_to_pes_6_sig_stat2trans(PENetwork_35_io_to_pes_6_sig_stat2trans),
    .io_to_pes_6_in_ready(PENetwork_35_io_to_pes_6_in_ready),
    .io_to_pes_6_out_ready(PENetwork_35_io_to_pes_6_out_ready),
    .io_to_pes_7_in_valid(PENetwork_35_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_35_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_35_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_35_io_to_pes_7_out_bits),
    .io_to_pes_7_sig_stat2trans(PENetwork_35_io_to_pes_7_sig_stat2trans),
    .io_to_pes_7_in_ready(PENetwork_35_io_to_pes_7_in_ready),
    .io_to_pes_7_out_ready(PENetwork_35_io_to_pes_7_out_ready),
    .io_to_pes_8_in_valid(PENetwork_35_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_35_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_35_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_35_io_to_pes_8_out_bits),
    .io_to_pes_8_sig_stat2trans(PENetwork_35_io_to_pes_8_sig_stat2trans),
    .io_to_pes_8_in_ready(PENetwork_35_io_to_pes_8_in_ready),
    .io_to_pes_8_out_ready(PENetwork_35_io_to_pes_8_out_ready),
    .io_to_pes_9_in_valid(PENetwork_35_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_35_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_35_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_35_io_to_pes_9_out_bits),
    .io_to_pes_9_sig_stat2trans(PENetwork_35_io_to_pes_9_sig_stat2trans),
    .io_to_pes_9_in_ready(PENetwork_35_io_to_pes_9_in_ready),
    .io_to_pes_9_out_ready(PENetwork_35_io_to_pes_9_out_ready),
    .io_to_pes_10_in_valid(PENetwork_35_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_35_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_35_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_35_io_to_pes_10_out_bits),
    .io_to_pes_10_sig_stat2trans(PENetwork_35_io_to_pes_10_sig_stat2trans),
    .io_to_pes_10_in_ready(PENetwork_35_io_to_pes_10_in_ready),
    .io_to_mem_valid(PENetwork_35_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_35_io_to_mem_bits),
    .io_sig_stat2trans(PENetwork_35_io_sig_stat2trans)
  );
  PENetwork_26 PENetwork_36 ( // @[pe.scala 227:13]
    .clock(PENetwork_36_clock),
    .io_to_pes_0_out_valid(PENetwork_36_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_36_io_to_pes_0_out_bits),
    .io_to_pes_0_sig_stat2trans(PENetwork_36_io_to_pes_0_sig_stat2trans),
    .io_to_pes_0_out_ready(PENetwork_36_io_to_pes_0_out_ready),
    .io_to_pes_1_in_valid(PENetwork_36_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_36_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_36_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_36_io_to_pes_1_out_bits),
    .io_to_pes_1_sig_stat2trans(PENetwork_36_io_to_pes_1_sig_stat2trans),
    .io_to_pes_1_in_ready(PENetwork_36_io_to_pes_1_in_ready),
    .io_to_pes_1_out_ready(PENetwork_36_io_to_pes_1_out_ready),
    .io_to_pes_2_in_valid(PENetwork_36_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_36_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_36_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_36_io_to_pes_2_out_bits),
    .io_to_pes_2_sig_stat2trans(PENetwork_36_io_to_pes_2_sig_stat2trans),
    .io_to_pes_2_in_ready(PENetwork_36_io_to_pes_2_in_ready),
    .io_to_pes_2_out_ready(PENetwork_36_io_to_pes_2_out_ready),
    .io_to_pes_3_in_valid(PENetwork_36_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_36_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_36_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_36_io_to_pes_3_out_bits),
    .io_to_pes_3_sig_stat2trans(PENetwork_36_io_to_pes_3_sig_stat2trans),
    .io_to_pes_3_in_ready(PENetwork_36_io_to_pes_3_in_ready),
    .io_to_pes_3_out_ready(PENetwork_36_io_to_pes_3_out_ready),
    .io_to_pes_4_in_valid(PENetwork_36_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_36_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_36_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_36_io_to_pes_4_out_bits),
    .io_to_pes_4_sig_stat2trans(PENetwork_36_io_to_pes_4_sig_stat2trans),
    .io_to_pes_4_in_ready(PENetwork_36_io_to_pes_4_in_ready),
    .io_to_pes_4_out_ready(PENetwork_36_io_to_pes_4_out_ready),
    .io_to_pes_5_in_valid(PENetwork_36_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_36_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_36_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_36_io_to_pes_5_out_bits),
    .io_to_pes_5_sig_stat2trans(PENetwork_36_io_to_pes_5_sig_stat2trans),
    .io_to_pes_5_in_ready(PENetwork_36_io_to_pes_5_in_ready),
    .io_to_pes_5_out_ready(PENetwork_36_io_to_pes_5_out_ready),
    .io_to_pes_6_in_valid(PENetwork_36_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_36_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_36_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_36_io_to_pes_6_out_bits),
    .io_to_pes_6_sig_stat2trans(PENetwork_36_io_to_pes_6_sig_stat2trans),
    .io_to_pes_6_in_ready(PENetwork_36_io_to_pes_6_in_ready),
    .io_to_pes_6_out_ready(PENetwork_36_io_to_pes_6_out_ready),
    .io_to_pes_7_in_valid(PENetwork_36_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_36_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_36_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_36_io_to_pes_7_out_bits),
    .io_to_pes_7_sig_stat2trans(PENetwork_36_io_to_pes_7_sig_stat2trans),
    .io_to_pes_7_in_ready(PENetwork_36_io_to_pes_7_in_ready),
    .io_to_pes_7_out_ready(PENetwork_36_io_to_pes_7_out_ready),
    .io_to_pes_8_in_valid(PENetwork_36_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_36_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_36_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_36_io_to_pes_8_out_bits),
    .io_to_pes_8_sig_stat2trans(PENetwork_36_io_to_pes_8_sig_stat2trans),
    .io_to_pes_8_in_ready(PENetwork_36_io_to_pes_8_in_ready),
    .io_to_pes_8_out_ready(PENetwork_36_io_to_pes_8_out_ready),
    .io_to_pes_9_in_valid(PENetwork_36_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_36_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_36_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_36_io_to_pes_9_out_bits),
    .io_to_pes_9_sig_stat2trans(PENetwork_36_io_to_pes_9_sig_stat2trans),
    .io_to_pes_9_in_ready(PENetwork_36_io_to_pes_9_in_ready),
    .io_to_pes_9_out_ready(PENetwork_36_io_to_pes_9_out_ready),
    .io_to_pes_10_in_valid(PENetwork_36_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_36_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_36_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_36_io_to_pes_10_out_bits),
    .io_to_pes_10_sig_stat2trans(PENetwork_36_io_to_pes_10_sig_stat2trans),
    .io_to_pes_10_in_ready(PENetwork_36_io_to_pes_10_in_ready),
    .io_to_mem_valid(PENetwork_36_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_36_io_to_mem_bits),
    .io_sig_stat2trans(PENetwork_36_io_sig_stat2trans)
  );
  PENetwork_26 PENetwork_37 ( // @[pe.scala 227:13]
    .clock(PENetwork_37_clock),
    .io_to_pes_0_out_valid(PENetwork_37_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_37_io_to_pes_0_out_bits),
    .io_to_pes_0_sig_stat2trans(PENetwork_37_io_to_pes_0_sig_stat2trans),
    .io_to_pes_0_out_ready(PENetwork_37_io_to_pes_0_out_ready),
    .io_to_pes_1_in_valid(PENetwork_37_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_37_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_37_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_37_io_to_pes_1_out_bits),
    .io_to_pes_1_sig_stat2trans(PENetwork_37_io_to_pes_1_sig_stat2trans),
    .io_to_pes_1_in_ready(PENetwork_37_io_to_pes_1_in_ready),
    .io_to_pes_1_out_ready(PENetwork_37_io_to_pes_1_out_ready),
    .io_to_pes_2_in_valid(PENetwork_37_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_37_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_37_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_37_io_to_pes_2_out_bits),
    .io_to_pes_2_sig_stat2trans(PENetwork_37_io_to_pes_2_sig_stat2trans),
    .io_to_pes_2_in_ready(PENetwork_37_io_to_pes_2_in_ready),
    .io_to_pes_2_out_ready(PENetwork_37_io_to_pes_2_out_ready),
    .io_to_pes_3_in_valid(PENetwork_37_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_37_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_37_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_37_io_to_pes_3_out_bits),
    .io_to_pes_3_sig_stat2trans(PENetwork_37_io_to_pes_3_sig_stat2trans),
    .io_to_pes_3_in_ready(PENetwork_37_io_to_pes_3_in_ready),
    .io_to_pes_3_out_ready(PENetwork_37_io_to_pes_3_out_ready),
    .io_to_pes_4_in_valid(PENetwork_37_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_37_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_37_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_37_io_to_pes_4_out_bits),
    .io_to_pes_4_sig_stat2trans(PENetwork_37_io_to_pes_4_sig_stat2trans),
    .io_to_pes_4_in_ready(PENetwork_37_io_to_pes_4_in_ready),
    .io_to_pes_4_out_ready(PENetwork_37_io_to_pes_4_out_ready),
    .io_to_pes_5_in_valid(PENetwork_37_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_37_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_37_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_37_io_to_pes_5_out_bits),
    .io_to_pes_5_sig_stat2trans(PENetwork_37_io_to_pes_5_sig_stat2trans),
    .io_to_pes_5_in_ready(PENetwork_37_io_to_pes_5_in_ready),
    .io_to_pes_5_out_ready(PENetwork_37_io_to_pes_5_out_ready),
    .io_to_pes_6_in_valid(PENetwork_37_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_37_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_37_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_37_io_to_pes_6_out_bits),
    .io_to_pes_6_sig_stat2trans(PENetwork_37_io_to_pes_6_sig_stat2trans),
    .io_to_pes_6_in_ready(PENetwork_37_io_to_pes_6_in_ready),
    .io_to_pes_6_out_ready(PENetwork_37_io_to_pes_6_out_ready),
    .io_to_pes_7_in_valid(PENetwork_37_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_37_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_37_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_37_io_to_pes_7_out_bits),
    .io_to_pes_7_sig_stat2trans(PENetwork_37_io_to_pes_7_sig_stat2trans),
    .io_to_pes_7_in_ready(PENetwork_37_io_to_pes_7_in_ready),
    .io_to_pes_7_out_ready(PENetwork_37_io_to_pes_7_out_ready),
    .io_to_pes_8_in_valid(PENetwork_37_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_37_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_37_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_37_io_to_pes_8_out_bits),
    .io_to_pes_8_sig_stat2trans(PENetwork_37_io_to_pes_8_sig_stat2trans),
    .io_to_pes_8_in_ready(PENetwork_37_io_to_pes_8_in_ready),
    .io_to_pes_8_out_ready(PENetwork_37_io_to_pes_8_out_ready),
    .io_to_pes_9_in_valid(PENetwork_37_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_37_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_37_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_37_io_to_pes_9_out_bits),
    .io_to_pes_9_sig_stat2trans(PENetwork_37_io_to_pes_9_sig_stat2trans),
    .io_to_pes_9_in_ready(PENetwork_37_io_to_pes_9_in_ready),
    .io_to_pes_9_out_ready(PENetwork_37_io_to_pes_9_out_ready),
    .io_to_pes_10_in_valid(PENetwork_37_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_37_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_37_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_37_io_to_pes_10_out_bits),
    .io_to_pes_10_sig_stat2trans(PENetwork_37_io_to_pes_10_sig_stat2trans),
    .io_to_pes_10_in_ready(PENetwork_37_io_to_pes_10_in_ready),
    .io_to_mem_valid(PENetwork_37_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_37_io_to_mem_bits),
    .io_sig_stat2trans(PENetwork_37_io_sig_stat2trans)
  );
  PENetwork_26 PENetwork_38 ( // @[pe.scala 227:13]
    .clock(PENetwork_38_clock),
    .io_to_pes_0_out_valid(PENetwork_38_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_38_io_to_pes_0_out_bits),
    .io_to_pes_0_sig_stat2trans(PENetwork_38_io_to_pes_0_sig_stat2trans),
    .io_to_pes_0_out_ready(PENetwork_38_io_to_pes_0_out_ready),
    .io_to_pes_1_in_valid(PENetwork_38_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_38_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_38_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_38_io_to_pes_1_out_bits),
    .io_to_pes_1_sig_stat2trans(PENetwork_38_io_to_pes_1_sig_stat2trans),
    .io_to_pes_1_in_ready(PENetwork_38_io_to_pes_1_in_ready),
    .io_to_pes_1_out_ready(PENetwork_38_io_to_pes_1_out_ready),
    .io_to_pes_2_in_valid(PENetwork_38_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_38_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_38_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_38_io_to_pes_2_out_bits),
    .io_to_pes_2_sig_stat2trans(PENetwork_38_io_to_pes_2_sig_stat2trans),
    .io_to_pes_2_in_ready(PENetwork_38_io_to_pes_2_in_ready),
    .io_to_pes_2_out_ready(PENetwork_38_io_to_pes_2_out_ready),
    .io_to_pes_3_in_valid(PENetwork_38_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_38_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_38_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_38_io_to_pes_3_out_bits),
    .io_to_pes_3_sig_stat2trans(PENetwork_38_io_to_pes_3_sig_stat2trans),
    .io_to_pes_3_in_ready(PENetwork_38_io_to_pes_3_in_ready),
    .io_to_pes_3_out_ready(PENetwork_38_io_to_pes_3_out_ready),
    .io_to_pes_4_in_valid(PENetwork_38_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_38_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_38_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_38_io_to_pes_4_out_bits),
    .io_to_pes_4_sig_stat2trans(PENetwork_38_io_to_pes_4_sig_stat2trans),
    .io_to_pes_4_in_ready(PENetwork_38_io_to_pes_4_in_ready),
    .io_to_pes_4_out_ready(PENetwork_38_io_to_pes_4_out_ready),
    .io_to_pes_5_in_valid(PENetwork_38_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_38_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_38_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_38_io_to_pes_5_out_bits),
    .io_to_pes_5_sig_stat2trans(PENetwork_38_io_to_pes_5_sig_stat2trans),
    .io_to_pes_5_in_ready(PENetwork_38_io_to_pes_5_in_ready),
    .io_to_pes_5_out_ready(PENetwork_38_io_to_pes_5_out_ready),
    .io_to_pes_6_in_valid(PENetwork_38_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_38_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_38_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_38_io_to_pes_6_out_bits),
    .io_to_pes_6_sig_stat2trans(PENetwork_38_io_to_pes_6_sig_stat2trans),
    .io_to_pes_6_in_ready(PENetwork_38_io_to_pes_6_in_ready),
    .io_to_pes_6_out_ready(PENetwork_38_io_to_pes_6_out_ready),
    .io_to_pes_7_in_valid(PENetwork_38_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_38_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_38_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_38_io_to_pes_7_out_bits),
    .io_to_pes_7_sig_stat2trans(PENetwork_38_io_to_pes_7_sig_stat2trans),
    .io_to_pes_7_in_ready(PENetwork_38_io_to_pes_7_in_ready),
    .io_to_pes_7_out_ready(PENetwork_38_io_to_pes_7_out_ready),
    .io_to_pes_8_in_valid(PENetwork_38_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_38_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_38_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_38_io_to_pes_8_out_bits),
    .io_to_pes_8_sig_stat2trans(PENetwork_38_io_to_pes_8_sig_stat2trans),
    .io_to_pes_8_in_ready(PENetwork_38_io_to_pes_8_in_ready),
    .io_to_pes_8_out_ready(PENetwork_38_io_to_pes_8_out_ready),
    .io_to_pes_9_in_valid(PENetwork_38_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_38_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_38_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_38_io_to_pes_9_out_bits),
    .io_to_pes_9_sig_stat2trans(PENetwork_38_io_to_pes_9_sig_stat2trans),
    .io_to_pes_9_in_ready(PENetwork_38_io_to_pes_9_in_ready),
    .io_to_pes_9_out_ready(PENetwork_38_io_to_pes_9_out_ready),
    .io_to_pes_10_in_valid(PENetwork_38_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_38_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_38_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_38_io_to_pes_10_out_bits),
    .io_to_pes_10_sig_stat2trans(PENetwork_38_io_to_pes_10_sig_stat2trans),
    .io_to_pes_10_in_ready(PENetwork_38_io_to_pes_10_in_ready),
    .io_to_mem_valid(PENetwork_38_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_38_io_to_mem_bits),
    .io_sig_stat2trans(PENetwork_38_io_sig_stat2trans)
  );
  PENetwork_26 PENetwork_39 ( // @[pe.scala 227:13]
    .clock(PENetwork_39_clock),
    .io_to_pes_0_out_valid(PENetwork_39_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_39_io_to_pes_0_out_bits),
    .io_to_pes_0_sig_stat2trans(PENetwork_39_io_to_pes_0_sig_stat2trans),
    .io_to_pes_0_out_ready(PENetwork_39_io_to_pes_0_out_ready),
    .io_to_pes_1_in_valid(PENetwork_39_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_39_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_39_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_39_io_to_pes_1_out_bits),
    .io_to_pes_1_sig_stat2trans(PENetwork_39_io_to_pes_1_sig_stat2trans),
    .io_to_pes_1_in_ready(PENetwork_39_io_to_pes_1_in_ready),
    .io_to_pes_1_out_ready(PENetwork_39_io_to_pes_1_out_ready),
    .io_to_pes_2_in_valid(PENetwork_39_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_39_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_39_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_39_io_to_pes_2_out_bits),
    .io_to_pes_2_sig_stat2trans(PENetwork_39_io_to_pes_2_sig_stat2trans),
    .io_to_pes_2_in_ready(PENetwork_39_io_to_pes_2_in_ready),
    .io_to_pes_2_out_ready(PENetwork_39_io_to_pes_2_out_ready),
    .io_to_pes_3_in_valid(PENetwork_39_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_39_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_39_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_39_io_to_pes_3_out_bits),
    .io_to_pes_3_sig_stat2trans(PENetwork_39_io_to_pes_3_sig_stat2trans),
    .io_to_pes_3_in_ready(PENetwork_39_io_to_pes_3_in_ready),
    .io_to_pes_3_out_ready(PENetwork_39_io_to_pes_3_out_ready),
    .io_to_pes_4_in_valid(PENetwork_39_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_39_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_39_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_39_io_to_pes_4_out_bits),
    .io_to_pes_4_sig_stat2trans(PENetwork_39_io_to_pes_4_sig_stat2trans),
    .io_to_pes_4_in_ready(PENetwork_39_io_to_pes_4_in_ready),
    .io_to_pes_4_out_ready(PENetwork_39_io_to_pes_4_out_ready),
    .io_to_pes_5_in_valid(PENetwork_39_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_39_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_39_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_39_io_to_pes_5_out_bits),
    .io_to_pes_5_sig_stat2trans(PENetwork_39_io_to_pes_5_sig_stat2trans),
    .io_to_pes_5_in_ready(PENetwork_39_io_to_pes_5_in_ready),
    .io_to_pes_5_out_ready(PENetwork_39_io_to_pes_5_out_ready),
    .io_to_pes_6_in_valid(PENetwork_39_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_39_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_39_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_39_io_to_pes_6_out_bits),
    .io_to_pes_6_sig_stat2trans(PENetwork_39_io_to_pes_6_sig_stat2trans),
    .io_to_pes_6_in_ready(PENetwork_39_io_to_pes_6_in_ready),
    .io_to_pes_6_out_ready(PENetwork_39_io_to_pes_6_out_ready),
    .io_to_pes_7_in_valid(PENetwork_39_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_39_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_39_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_39_io_to_pes_7_out_bits),
    .io_to_pes_7_sig_stat2trans(PENetwork_39_io_to_pes_7_sig_stat2trans),
    .io_to_pes_7_in_ready(PENetwork_39_io_to_pes_7_in_ready),
    .io_to_pes_7_out_ready(PENetwork_39_io_to_pes_7_out_ready),
    .io_to_pes_8_in_valid(PENetwork_39_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_39_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_39_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_39_io_to_pes_8_out_bits),
    .io_to_pes_8_sig_stat2trans(PENetwork_39_io_to_pes_8_sig_stat2trans),
    .io_to_pes_8_in_ready(PENetwork_39_io_to_pes_8_in_ready),
    .io_to_pes_8_out_ready(PENetwork_39_io_to_pes_8_out_ready),
    .io_to_pes_9_in_valid(PENetwork_39_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_39_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_39_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_39_io_to_pes_9_out_bits),
    .io_to_pes_9_sig_stat2trans(PENetwork_39_io_to_pes_9_sig_stat2trans),
    .io_to_pes_9_in_ready(PENetwork_39_io_to_pes_9_in_ready),
    .io_to_pes_9_out_ready(PENetwork_39_io_to_pes_9_out_ready),
    .io_to_pes_10_in_valid(PENetwork_39_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_39_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_39_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_39_io_to_pes_10_out_bits),
    .io_to_pes_10_sig_stat2trans(PENetwork_39_io_to_pes_10_sig_stat2trans),
    .io_to_pes_10_in_ready(PENetwork_39_io_to_pes_10_in_ready),
    .io_to_mem_valid(PENetwork_39_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_39_io_to_mem_bits),
    .io_sig_stat2trans(PENetwork_39_io_sig_stat2trans)
  );
  PENetwork_26 PENetwork_40 ( // @[pe.scala 227:13]
    .clock(PENetwork_40_clock),
    .io_to_pes_0_out_valid(PENetwork_40_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_40_io_to_pes_0_out_bits),
    .io_to_pes_0_sig_stat2trans(PENetwork_40_io_to_pes_0_sig_stat2trans),
    .io_to_pes_0_out_ready(PENetwork_40_io_to_pes_0_out_ready),
    .io_to_pes_1_in_valid(PENetwork_40_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_40_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_40_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_40_io_to_pes_1_out_bits),
    .io_to_pes_1_sig_stat2trans(PENetwork_40_io_to_pes_1_sig_stat2trans),
    .io_to_pes_1_in_ready(PENetwork_40_io_to_pes_1_in_ready),
    .io_to_pes_1_out_ready(PENetwork_40_io_to_pes_1_out_ready),
    .io_to_pes_2_in_valid(PENetwork_40_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_40_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_40_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_40_io_to_pes_2_out_bits),
    .io_to_pes_2_sig_stat2trans(PENetwork_40_io_to_pes_2_sig_stat2trans),
    .io_to_pes_2_in_ready(PENetwork_40_io_to_pes_2_in_ready),
    .io_to_pes_2_out_ready(PENetwork_40_io_to_pes_2_out_ready),
    .io_to_pes_3_in_valid(PENetwork_40_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_40_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_40_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_40_io_to_pes_3_out_bits),
    .io_to_pes_3_sig_stat2trans(PENetwork_40_io_to_pes_3_sig_stat2trans),
    .io_to_pes_3_in_ready(PENetwork_40_io_to_pes_3_in_ready),
    .io_to_pes_3_out_ready(PENetwork_40_io_to_pes_3_out_ready),
    .io_to_pes_4_in_valid(PENetwork_40_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_40_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_40_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_40_io_to_pes_4_out_bits),
    .io_to_pes_4_sig_stat2trans(PENetwork_40_io_to_pes_4_sig_stat2trans),
    .io_to_pes_4_in_ready(PENetwork_40_io_to_pes_4_in_ready),
    .io_to_pes_4_out_ready(PENetwork_40_io_to_pes_4_out_ready),
    .io_to_pes_5_in_valid(PENetwork_40_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_40_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_40_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_40_io_to_pes_5_out_bits),
    .io_to_pes_5_sig_stat2trans(PENetwork_40_io_to_pes_5_sig_stat2trans),
    .io_to_pes_5_in_ready(PENetwork_40_io_to_pes_5_in_ready),
    .io_to_pes_5_out_ready(PENetwork_40_io_to_pes_5_out_ready),
    .io_to_pes_6_in_valid(PENetwork_40_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_40_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_40_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_40_io_to_pes_6_out_bits),
    .io_to_pes_6_sig_stat2trans(PENetwork_40_io_to_pes_6_sig_stat2trans),
    .io_to_pes_6_in_ready(PENetwork_40_io_to_pes_6_in_ready),
    .io_to_pes_6_out_ready(PENetwork_40_io_to_pes_6_out_ready),
    .io_to_pes_7_in_valid(PENetwork_40_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_40_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_40_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_40_io_to_pes_7_out_bits),
    .io_to_pes_7_sig_stat2trans(PENetwork_40_io_to_pes_7_sig_stat2trans),
    .io_to_pes_7_in_ready(PENetwork_40_io_to_pes_7_in_ready),
    .io_to_pes_7_out_ready(PENetwork_40_io_to_pes_7_out_ready),
    .io_to_pes_8_in_valid(PENetwork_40_io_to_pes_8_in_valid),
    .io_to_pes_8_in_bits(PENetwork_40_io_to_pes_8_in_bits),
    .io_to_pes_8_out_valid(PENetwork_40_io_to_pes_8_out_valid),
    .io_to_pes_8_out_bits(PENetwork_40_io_to_pes_8_out_bits),
    .io_to_pes_8_sig_stat2trans(PENetwork_40_io_to_pes_8_sig_stat2trans),
    .io_to_pes_8_in_ready(PENetwork_40_io_to_pes_8_in_ready),
    .io_to_pes_8_out_ready(PENetwork_40_io_to_pes_8_out_ready),
    .io_to_pes_9_in_valid(PENetwork_40_io_to_pes_9_in_valid),
    .io_to_pes_9_in_bits(PENetwork_40_io_to_pes_9_in_bits),
    .io_to_pes_9_out_valid(PENetwork_40_io_to_pes_9_out_valid),
    .io_to_pes_9_out_bits(PENetwork_40_io_to_pes_9_out_bits),
    .io_to_pes_9_sig_stat2trans(PENetwork_40_io_to_pes_9_sig_stat2trans),
    .io_to_pes_9_in_ready(PENetwork_40_io_to_pes_9_in_ready),
    .io_to_pes_9_out_ready(PENetwork_40_io_to_pes_9_out_ready),
    .io_to_pes_10_in_valid(PENetwork_40_io_to_pes_10_in_valid),
    .io_to_pes_10_in_bits(PENetwork_40_io_to_pes_10_in_bits),
    .io_to_pes_10_out_valid(PENetwork_40_io_to_pes_10_out_valid),
    .io_to_pes_10_out_bits(PENetwork_40_io_to_pes_10_out_bits),
    .io_to_pes_10_sig_stat2trans(PENetwork_40_io_to_pes_10_sig_stat2trans),
    .io_to_pes_10_in_ready(PENetwork_40_io_to_pes_10_in_ready),
    .io_to_mem_valid(PENetwork_40_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_40_io_to_mem_bits),
    .io_sig_stat2trans(PENetwork_40_io_sig_stat2trans)
  );
  MemController MemController ( // @[pe.scala 306:15]
    .clock(MemController_clock),
    .reset(MemController_reset),
    .io_rd_valid(MemController_io_rd_valid),
    .io_wr_valid(MemController_io_wr_valid),
    .io_rd_data_valid(MemController_io_rd_data_valid),
    .io_rd_data_bits(MemController_io_rd_data_bits),
    .io_wr_data_valid(MemController_io_wr_data_valid),
    .io_wr_data_bits(MemController_io_wr_data_bits)
  );
  MemController MemController_1 ( // @[pe.scala 306:15]
    .clock(MemController_1_clock),
    .reset(MemController_1_reset),
    .io_rd_valid(MemController_1_io_rd_valid),
    .io_wr_valid(MemController_1_io_wr_valid),
    .io_rd_data_valid(MemController_1_io_rd_data_valid),
    .io_rd_data_bits(MemController_1_io_rd_data_bits),
    .io_wr_data_valid(MemController_1_io_wr_data_valid),
    .io_wr_data_bits(MemController_1_io_wr_data_bits)
  );
  MemController MemController_2 ( // @[pe.scala 306:15]
    .clock(MemController_2_clock),
    .reset(MemController_2_reset),
    .io_rd_valid(MemController_2_io_rd_valid),
    .io_wr_valid(MemController_2_io_wr_valid),
    .io_rd_data_valid(MemController_2_io_rd_data_valid),
    .io_rd_data_bits(MemController_2_io_rd_data_bits),
    .io_wr_data_valid(MemController_2_io_wr_data_valid),
    .io_wr_data_bits(MemController_2_io_wr_data_bits)
  );
  MemController MemController_3 ( // @[pe.scala 306:15]
    .clock(MemController_3_clock),
    .reset(MemController_3_reset),
    .io_rd_valid(MemController_3_io_rd_valid),
    .io_wr_valid(MemController_3_io_wr_valid),
    .io_rd_data_valid(MemController_3_io_rd_data_valid),
    .io_rd_data_bits(MemController_3_io_rd_data_bits),
    .io_wr_data_valid(MemController_3_io_wr_data_valid),
    .io_wr_data_bits(MemController_3_io_wr_data_bits)
  );
  MemController MemController_4 ( // @[pe.scala 306:15]
    .clock(MemController_4_clock),
    .reset(MemController_4_reset),
    .io_rd_valid(MemController_4_io_rd_valid),
    .io_wr_valid(MemController_4_io_wr_valid),
    .io_rd_data_valid(MemController_4_io_rd_data_valid),
    .io_rd_data_bits(MemController_4_io_rd_data_bits),
    .io_wr_data_valid(MemController_4_io_wr_data_valid),
    .io_wr_data_bits(MemController_4_io_wr_data_bits)
  );
  MemController MemController_5 ( // @[pe.scala 306:15]
    .clock(MemController_5_clock),
    .reset(MemController_5_reset),
    .io_rd_valid(MemController_5_io_rd_valid),
    .io_wr_valid(MemController_5_io_wr_valid),
    .io_rd_data_valid(MemController_5_io_rd_data_valid),
    .io_rd_data_bits(MemController_5_io_rd_data_bits),
    .io_wr_data_valid(MemController_5_io_wr_data_valid),
    .io_wr_data_bits(MemController_5_io_wr_data_bits)
  );
  MemController MemController_6 ( // @[pe.scala 306:15]
    .clock(MemController_6_clock),
    .reset(MemController_6_reset),
    .io_rd_valid(MemController_6_io_rd_valid),
    .io_wr_valid(MemController_6_io_wr_valid),
    .io_rd_data_valid(MemController_6_io_rd_data_valid),
    .io_rd_data_bits(MemController_6_io_rd_data_bits),
    .io_wr_data_valid(MemController_6_io_wr_data_valid),
    .io_wr_data_bits(MemController_6_io_wr_data_bits)
  );
  MemController MemController_7 ( // @[pe.scala 306:15]
    .clock(MemController_7_clock),
    .reset(MemController_7_reset),
    .io_rd_valid(MemController_7_io_rd_valid),
    .io_wr_valid(MemController_7_io_wr_valid),
    .io_rd_data_valid(MemController_7_io_rd_data_valid),
    .io_rd_data_bits(MemController_7_io_rd_data_bits),
    .io_wr_data_valid(MemController_7_io_wr_data_valid),
    .io_wr_data_bits(MemController_7_io_wr_data_bits)
  );
  MemController MemController_8 ( // @[pe.scala 306:15]
    .clock(MemController_8_clock),
    .reset(MemController_8_reset),
    .io_rd_valid(MemController_8_io_rd_valid),
    .io_wr_valid(MemController_8_io_wr_valid),
    .io_rd_data_valid(MemController_8_io_rd_data_valid),
    .io_rd_data_bits(MemController_8_io_rd_data_bits),
    .io_wr_data_valid(MemController_8_io_wr_data_valid),
    .io_wr_data_bits(MemController_8_io_wr_data_bits)
  );
  MemController MemController_9 ( // @[pe.scala 306:15]
    .clock(MemController_9_clock),
    .reset(MemController_9_reset),
    .io_rd_valid(MemController_9_io_rd_valid),
    .io_wr_valid(MemController_9_io_wr_valid),
    .io_rd_data_valid(MemController_9_io_rd_data_valid),
    .io_rd_data_bits(MemController_9_io_rd_data_bits),
    .io_wr_data_valid(MemController_9_io_wr_data_valid),
    .io_wr_data_bits(MemController_9_io_wr_data_bits)
  );
  MemController MemController_10 ( // @[pe.scala 306:15]
    .clock(MemController_10_clock),
    .reset(MemController_10_reset),
    .io_rd_valid(MemController_10_io_rd_valid),
    .io_wr_valid(MemController_10_io_wr_valid),
    .io_rd_data_valid(MemController_10_io_rd_data_valid),
    .io_rd_data_bits(MemController_10_io_rd_data_bits),
    .io_wr_data_valid(MemController_10_io_wr_data_valid),
    .io_wr_data_bits(MemController_10_io_wr_data_bits)
  );
  MemController_11 MemController_11 ( // @[pe.scala 306:15]
    .clock(MemController_11_clock),
    .reset(MemController_11_reset),
    .io_rd_valid(MemController_11_io_rd_valid),
    .io_wr_valid(MemController_11_io_wr_valid),
    .io_rd_data_valid(MemController_11_io_rd_data_valid),
    .io_rd_data_bits(MemController_11_io_rd_data_bits),
    .io_wr_data_valid(MemController_11_io_wr_data_valid),
    .io_wr_data_bits(MemController_11_io_wr_data_bits)
  );
  MemController_11 MemController_12 ( // @[pe.scala 306:15]
    .clock(MemController_12_clock),
    .reset(MemController_12_reset),
    .io_rd_valid(MemController_12_io_rd_valid),
    .io_wr_valid(MemController_12_io_wr_valid),
    .io_rd_data_valid(MemController_12_io_rd_data_valid),
    .io_rd_data_bits(MemController_12_io_rd_data_bits),
    .io_wr_data_valid(MemController_12_io_wr_data_valid),
    .io_wr_data_bits(MemController_12_io_wr_data_bits)
  );
  MemController_11 MemController_13 ( // @[pe.scala 306:15]
    .clock(MemController_13_clock),
    .reset(MemController_13_reset),
    .io_rd_valid(MemController_13_io_rd_valid),
    .io_wr_valid(MemController_13_io_wr_valid),
    .io_rd_data_valid(MemController_13_io_rd_data_valid),
    .io_rd_data_bits(MemController_13_io_rd_data_bits),
    .io_wr_data_valid(MemController_13_io_wr_data_valid),
    .io_wr_data_bits(MemController_13_io_wr_data_bits)
  );
  MemController_11 MemController_14 ( // @[pe.scala 306:15]
    .clock(MemController_14_clock),
    .reset(MemController_14_reset),
    .io_rd_valid(MemController_14_io_rd_valid),
    .io_wr_valid(MemController_14_io_wr_valid),
    .io_rd_data_valid(MemController_14_io_rd_data_valid),
    .io_rd_data_bits(MemController_14_io_rd_data_bits),
    .io_wr_data_valid(MemController_14_io_wr_data_valid),
    .io_wr_data_bits(MemController_14_io_wr_data_bits)
  );
  MemController_11 MemController_15 ( // @[pe.scala 306:15]
    .clock(MemController_15_clock),
    .reset(MemController_15_reset),
    .io_rd_valid(MemController_15_io_rd_valid),
    .io_wr_valid(MemController_15_io_wr_valid),
    .io_rd_data_valid(MemController_15_io_rd_data_valid),
    .io_rd_data_bits(MemController_15_io_rd_data_bits),
    .io_wr_data_valid(MemController_15_io_wr_data_valid),
    .io_wr_data_bits(MemController_15_io_wr_data_bits)
  );
  MemController_11 MemController_16 ( // @[pe.scala 306:15]
    .clock(MemController_16_clock),
    .reset(MemController_16_reset),
    .io_rd_valid(MemController_16_io_rd_valid),
    .io_wr_valid(MemController_16_io_wr_valid),
    .io_rd_data_valid(MemController_16_io_rd_data_valid),
    .io_rd_data_bits(MemController_16_io_rd_data_bits),
    .io_wr_data_valid(MemController_16_io_wr_data_valid),
    .io_wr_data_bits(MemController_16_io_wr_data_bits)
  );
  MemController_11 MemController_17 ( // @[pe.scala 306:15]
    .clock(MemController_17_clock),
    .reset(MemController_17_reset),
    .io_rd_valid(MemController_17_io_rd_valid),
    .io_wr_valid(MemController_17_io_wr_valid),
    .io_rd_data_valid(MemController_17_io_rd_data_valid),
    .io_rd_data_bits(MemController_17_io_rd_data_bits),
    .io_wr_data_valid(MemController_17_io_wr_data_valid),
    .io_wr_data_bits(MemController_17_io_wr_data_bits)
  );
  MemController_11 MemController_18 ( // @[pe.scala 306:15]
    .clock(MemController_18_clock),
    .reset(MemController_18_reset),
    .io_rd_valid(MemController_18_io_rd_valid),
    .io_wr_valid(MemController_18_io_wr_valid),
    .io_rd_data_valid(MemController_18_io_rd_data_valid),
    .io_rd_data_bits(MemController_18_io_rd_data_bits),
    .io_wr_data_valid(MemController_18_io_wr_data_valid),
    .io_wr_data_bits(MemController_18_io_wr_data_bits)
  );
  MemController_11 MemController_19 ( // @[pe.scala 306:15]
    .clock(MemController_19_clock),
    .reset(MemController_19_reset),
    .io_rd_valid(MemController_19_io_rd_valid),
    .io_wr_valid(MemController_19_io_wr_valid),
    .io_rd_data_valid(MemController_19_io_rd_data_valid),
    .io_rd_data_bits(MemController_19_io_rd_data_bits),
    .io_wr_data_valid(MemController_19_io_wr_data_valid),
    .io_wr_data_bits(MemController_19_io_wr_data_bits)
  );
  MemController_11 MemController_20 ( // @[pe.scala 306:15]
    .clock(MemController_20_clock),
    .reset(MemController_20_reset),
    .io_rd_valid(MemController_20_io_rd_valid),
    .io_wr_valid(MemController_20_io_wr_valid),
    .io_rd_data_valid(MemController_20_io_rd_data_valid),
    .io_rd_data_bits(MemController_20_io_rd_data_bits),
    .io_wr_data_valid(MemController_20_io_wr_data_valid),
    .io_wr_data_bits(MemController_20_io_wr_data_bits)
  );
  MemController_11 MemController_21 ( // @[pe.scala 306:15]
    .clock(MemController_21_clock),
    .reset(MemController_21_reset),
    .io_rd_valid(MemController_21_io_rd_valid),
    .io_wr_valid(MemController_21_io_wr_valid),
    .io_rd_data_valid(MemController_21_io_rd_data_valid),
    .io_rd_data_bits(MemController_21_io_rd_data_bits),
    .io_wr_data_valid(MemController_21_io_wr_data_valid),
    .io_wr_data_bits(MemController_21_io_wr_data_bits)
  );
  MemController_11 MemController_22 ( // @[pe.scala 306:15]
    .clock(MemController_22_clock),
    .reset(MemController_22_reset),
    .io_rd_valid(MemController_22_io_rd_valid),
    .io_wr_valid(MemController_22_io_wr_valid),
    .io_rd_data_valid(MemController_22_io_rd_data_valid),
    .io_rd_data_bits(MemController_22_io_rd_data_bits),
    .io_wr_data_valid(MemController_22_io_wr_data_valid),
    .io_wr_data_bits(MemController_22_io_wr_data_bits)
  );
  MemController_11 MemController_23 ( // @[pe.scala 306:15]
    .clock(MemController_23_clock),
    .reset(MemController_23_reset),
    .io_rd_valid(MemController_23_io_rd_valid),
    .io_wr_valid(MemController_23_io_wr_valid),
    .io_rd_data_valid(MemController_23_io_rd_data_valid),
    .io_rd_data_bits(MemController_23_io_rd_data_bits),
    .io_wr_data_valid(MemController_23_io_wr_data_valid),
    .io_wr_data_bits(MemController_23_io_wr_data_bits)
  );
  MemController_11 MemController_24 ( // @[pe.scala 306:15]
    .clock(MemController_24_clock),
    .reset(MemController_24_reset),
    .io_rd_valid(MemController_24_io_rd_valid),
    .io_wr_valid(MemController_24_io_wr_valid),
    .io_rd_data_valid(MemController_24_io_rd_data_valid),
    .io_rd_data_bits(MemController_24_io_rd_data_bits),
    .io_wr_data_valid(MemController_24_io_wr_data_valid),
    .io_wr_data_bits(MemController_24_io_wr_data_bits)
  );
  MemController_11 MemController_25 ( // @[pe.scala 306:15]
    .clock(MemController_25_clock),
    .reset(MemController_25_reset),
    .io_rd_valid(MemController_25_io_rd_valid),
    .io_wr_valid(MemController_25_io_wr_valid),
    .io_rd_data_valid(MemController_25_io_rd_data_valid),
    .io_rd_data_bits(MemController_25_io_rd_data_bits),
    .io_wr_data_valid(MemController_25_io_wr_data_valid),
    .io_wr_data_bits(MemController_25_io_wr_data_bits)
  );
  MemController_26 MemController_26 ( // @[pe.scala 304:15]
    .clock(MemController_26_clock),
    .reset(MemController_26_reset),
    .io_rd_valid(MemController_26_io_rd_valid),
    .io_wr_valid(MemController_26_io_wr_valid),
    .io_rd_data_valid(MemController_26_io_rd_data_valid),
    .io_rd_data_bits(MemController_26_io_rd_data_bits),
    .io_wr_data_valid(MemController_26_io_wr_data_valid),
    .io_wr_data_bits(MemController_26_io_wr_data_bits)
  );
  MemController_26 MemController_27 ( // @[pe.scala 304:15]
    .clock(MemController_27_clock),
    .reset(MemController_27_reset),
    .io_rd_valid(MemController_27_io_rd_valid),
    .io_wr_valid(MemController_27_io_wr_valid),
    .io_rd_data_valid(MemController_27_io_rd_data_valid),
    .io_rd_data_bits(MemController_27_io_rd_data_bits),
    .io_wr_data_valid(MemController_27_io_wr_data_valid),
    .io_wr_data_bits(MemController_27_io_wr_data_bits)
  );
  MemController_26 MemController_28 ( // @[pe.scala 304:15]
    .clock(MemController_28_clock),
    .reset(MemController_28_reset),
    .io_rd_valid(MemController_28_io_rd_valid),
    .io_wr_valid(MemController_28_io_wr_valid),
    .io_rd_data_valid(MemController_28_io_rd_data_valid),
    .io_rd_data_bits(MemController_28_io_rd_data_bits),
    .io_wr_data_valid(MemController_28_io_wr_data_valid),
    .io_wr_data_bits(MemController_28_io_wr_data_bits)
  );
  MemController_26 MemController_29 ( // @[pe.scala 304:15]
    .clock(MemController_29_clock),
    .reset(MemController_29_reset),
    .io_rd_valid(MemController_29_io_rd_valid),
    .io_wr_valid(MemController_29_io_wr_valid),
    .io_rd_data_valid(MemController_29_io_rd_data_valid),
    .io_rd_data_bits(MemController_29_io_rd_data_bits),
    .io_wr_data_valid(MemController_29_io_wr_data_valid),
    .io_wr_data_bits(MemController_29_io_wr_data_bits)
  );
  MemController_26 MemController_30 ( // @[pe.scala 304:15]
    .clock(MemController_30_clock),
    .reset(MemController_30_reset),
    .io_rd_valid(MemController_30_io_rd_valid),
    .io_wr_valid(MemController_30_io_wr_valid),
    .io_rd_data_valid(MemController_30_io_rd_data_valid),
    .io_rd_data_bits(MemController_30_io_rd_data_bits),
    .io_wr_data_valid(MemController_30_io_wr_data_valid),
    .io_wr_data_bits(MemController_30_io_wr_data_bits)
  );
  MemController_26 MemController_31 ( // @[pe.scala 304:15]
    .clock(MemController_31_clock),
    .reset(MemController_31_reset),
    .io_rd_valid(MemController_31_io_rd_valid),
    .io_wr_valid(MemController_31_io_wr_valid),
    .io_rd_data_valid(MemController_31_io_rd_data_valid),
    .io_rd_data_bits(MemController_31_io_rd_data_bits),
    .io_wr_data_valid(MemController_31_io_wr_data_valid),
    .io_wr_data_bits(MemController_31_io_wr_data_bits)
  );
  MemController_26 MemController_32 ( // @[pe.scala 304:15]
    .clock(MemController_32_clock),
    .reset(MemController_32_reset),
    .io_rd_valid(MemController_32_io_rd_valid),
    .io_wr_valid(MemController_32_io_wr_valid),
    .io_rd_data_valid(MemController_32_io_rd_data_valid),
    .io_rd_data_bits(MemController_32_io_rd_data_bits),
    .io_wr_data_valid(MemController_32_io_wr_data_valid),
    .io_wr_data_bits(MemController_32_io_wr_data_bits)
  );
  MemController_26 MemController_33 ( // @[pe.scala 304:15]
    .clock(MemController_33_clock),
    .reset(MemController_33_reset),
    .io_rd_valid(MemController_33_io_rd_valid),
    .io_wr_valid(MemController_33_io_wr_valid),
    .io_rd_data_valid(MemController_33_io_rd_data_valid),
    .io_rd_data_bits(MemController_33_io_rd_data_bits),
    .io_wr_data_valid(MemController_33_io_wr_data_valid),
    .io_wr_data_bits(MemController_33_io_wr_data_bits)
  );
  MemController_26 MemController_34 ( // @[pe.scala 304:15]
    .clock(MemController_34_clock),
    .reset(MemController_34_reset),
    .io_rd_valid(MemController_34_io_rd_valid),
    .io_wr_valid(MemController_34_io_wr_valid),
    .io_rd_data_valid(MemController_34_io_rd_data_valid),
    .io_rd_data_bits(MemController_34_io_rd_data_bits),
    .io_wr_data_valid(MemController_34_io_wr_data_valid),
    .io_wr_data_bits(MemController_34_io_wr_data_bits)
  );
  MemController_26 MemController_35 ( // @[pe.scala 304:15]
    .clock(MemController_35_clock),
    .reset(MemController_35_reset),
    .io_rd_valid(MemController_35_io_rd_valid),
    .io_wr_valid(MemController_35_io_wr_valid),
    .io_rd_data_valid(MemController_35_io_rd_data_valid),
    .io_rd_data_bits(MemController_35_io_rd_data_bits),
    .io_wr_data_valid(MemController_35_io_wr_data_valid),
    .io_wr_data_bits(MemController_35_io_wr_data_bits)
  );
  MemController_26 MemController_36 ( // @[pe.scala 304:15]
    .clock(MemController_36_clock),
    .reset(MemController_36_reset),
    .io_rd_valid(MemController_36_io_rd_valid),
    .io_wr_valid(MemController_36_io_wr_valid),
    .io_rd_data_valid(MemController_36_io_rd_data_valid),
    .io_rd_data_bits(MemController_36_io_rd_data_bits),
    .io_wr_data_valid(MemController_36_io_wr_data_valid),
    .io_wr_data_bits(MemController_36_io_wr_data_bits)
  );
  MemController_26 MemController_37 ( // @[pe.scala 304:15]
    .clock(MemController_37_clock),
    .reset(MemController_37_reset),
    .io_rd_valid(MemController_37_io_rd_valid),
    .io_wr_valid(MemController_37_io_wr_valid),
    .io_rd_data_valid(MemController_37_io_rd_data_valid),
    .io_rd_data_bits(MemController_37_io_rd_data_bits),
    .io_wr_data_valid(MemController_37_io_wr_data_valid),
    .io_wr_data_bits(MemController_37_io_wr_data_bits)
  );
  MemController_26 MemController_38 ( // @[pe.scala 304:15]
    .clock(MemController_38_clock),
    .reset(MemController_38_reset),
    .io_rd_valid(MemController_38_io_rd_valid),
    .io_wr_valid(MemController_38_io_wr_valid),
    .io_rd_data_valid(MemController_38_io_rd_data_valid),
    .io_rd_data_bits(MemController_38_io_rd_data_bits),
    .io_wr_data_valid(MemController_38_io_wr_data_valid),
    .io_wr_data_bits(MemController_38_io_wr_data_bits)
  );
  MemController_26 MemController_39 ( // @[pe.scala 304:15]
    .clock(MemController_39_clock),
    .reset(MemController_39_reset),
    .io_rd_valid(MemController_39_io_rd_valid),
    .io_wr_valid(MemController_39_io_wr_valid),
    .io_rd_data_valid(MemController_39_io_rd_data_valid),
    .io_rd_data_bits(MemController_39_io_rd_data_bits),
    .io_wr_data_valid(MemController_39_io_wr_data_valid),
    .io_wr_data_bits(MemController_39_io_wr_data_bits)
  );
  MemController_26 MemController_40 ( // @[pe.scala 304:15]
    .clock(MemController_40_clock),
    .reset(MemController_40_reset),
    .io_rd_valid(MemController_40_io_rd_valid),
    .io_wr_valid(MemController_40_io_wr_valid),
    .io_rd_data_valid(MemController_40_io_rd_data_valid),
    .io_rd_data_bits(MemController_40_io_rd_data_bits),
    .io_wr_data_valid(MemController_40_io_wr_data_valid),
    .io_wr_data_bits(MemController_40_io_wr_data_bits)
  );
  assign io_data_2_out_0_valid = MemController_26_io_rd_data_valid; // @[pe.scala 321:31]
  assign io_data_2_out_0_bits = MemController_26_io_rd_data_bits; // @[pe.scala 321:31]
  assign io_data_2_out_1_valid = MemController_27_io_rd_data_valid; // @[pe.scala 321:31]
  assign io_data_2_out_1_bits = MemController_27_io_rd_data_bits; // @[pe.scala 321:31]
  assign io_data_2_out_2_valid = MemController_28_io_rd_data_valid; // @[pe.scala 321:31]
  assign io_data_2_out_2_bits = MemController_28_io_rd_data_bits; // @[pe.scala 321:31]
  assign io_data_2_out_3_valid = MemController_29_io_rd_data_valid; // @[pe.scala 321:31]
  assign io_data_2_out_3_bits = MemController_29_io_rd_data_bits; // @[pe.scala 321:31]
  assign io_data_2_out_4_valid = MemController_30_io_rd_data_valid; // @[pe.scala 321:31]
  assign io_data_2_out_4_bits = MemController_30_io_rd_data_bits; // @[pe.scala 321:31]
  assign io_data_2_out_5_valid = MemController_31_io_rd_data_valid; // @[pe.scala 321:31]
  assign io_data_2_out_5_bits = MemController_31_io_rd_data_bits; // @[pe.scala 321:31]
  assign io_data_2_out_6_valid = MemController_32_io_rd_data_valid; // @[pe.scala 321:31]
  assign io_data_2_out_6_bits = MemController_32_io_rd_data_bits; // @[pe.scala 321:31]
  assign io_data_2_out_7_valid = MemController_33_io_rd_data_valid; // @[pe.scala 321:31]
  assign io_data_2_out_7_bits = MemController_33_io_rd_data_bits; // @[pe.scala 321:31]
  assign io_data_2_out_8_valid = MemController_34_io_rd_data_valid; // @[pe.scala 321:31]
  assign io_data_2_out_8_bits = MemController_34_io_rd_data_bits; // @[pe.scala 321:31]
  assign io_data_2_out_9_valid = MemController_35_io_rd_data_valid; // @[pe.scala 321:31]
  assign io_data_2_out_9_bits = MemController_35_io_rd_data_bits; // @[pe.scala 321:31]
  assign io_data_2_out_10_valid = MemController_36_io_rd_data_valid; // @[pe.scala 321:31]
  assign io_data_2_out_10_bits = MemController_36_io_rd_data_bits; // @[pe.scala 321:31]
  assign io_data_2_out_11_valid = MemController_37_io_rd_data_valid; // @[pe.scala 321:31]
  assign io_data_2_out_11_bits = MemController_37_io_rd_data_bits; // @[pe.scala 321:31]
  assign io_data_2_out_12_valid = MemController_38_io_rd_data_valid; // @[pe.scala 321:31]
  assign io_data_2_out_12_bits = MemController_38_io_rd_data_bits; // @[pe.scala 321:31]
  assign io_data_2_out_13_valid = MemController_39_io_rd_data_valid; // @[pe.scala 321:31]
  assign io_data_2_out_13_bits = MemController_39_io_rd_data_bits; // @[pe.scala 321:31]
  assign io_data_2_out_14_valid = MemController_40_io_rd_data_valid; // @[pe.scala 321:31]
  assign io_data_2_out_14_bits = MemController_40_io_rd_data_bits; // @[pe.scala 321:31]
  assign MultiDimTime_clock = clock;
  assign MultiDimTime_reset = reset;
  assign MultiDimTime_io_in = io_exec_valid; // @[pe.scala 255:16]
  assign PE_clock = clock;
  assign PE_reset = reset;
  assign PE_io_data_2_in_valid = 1'h0; // @[pe.scala 262:34]
  assign PE_io_data_2_in_bits = 256'h0; // @[pe.scala 262:34]
  assign PE_io_data_2_sig_stat2trans = PENetwork_26_io_to_pes_0_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_io_data_2_out_ready = PENetwork_26_io_to_pes_0_out_ready; // @[pe.scala 268:49]
  assign PE_io_data_1_in_valid = PENetwork_11_io_to_pes_0_in_valid; // @[pe.scala 262:34]
  assign PE_io_data_1_in_bits = PENetwork_11_io_to_pes_0_in_bits; // @[pe.scala 262:34]
  assign PE_io_data_0_in_valid = PENetwork_io_to_pes_0_in_valid; // @[pe.scala 262:34]
  assign PE_io_data_0_in_bits = PENetwork_io_to_pes_0_in_bits; // @[pe.scala 262:34]
  assign PE_1_clock = clock;
  assign PE_1_reset = reset;
  assign PE_1_io_data_2_in_valid = PENetwork_26_io_to_pes_1_in_valid; // @[pe.scala 262:34]
  assign PE_1_io_data_2_in_bits = PENetwork_26_io_to_pes_1_in_bits; // @[pe.scala 262:34]
  assign PE_1_io_data_2_sig_stat2trans = PENetwork_26_io_to_pes_1_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_1_io_data_2_out_ready = PENetwork_26_io_to_pes_1_out_ready; // @[pe.scala 268:49]
  assign PE_1_io_data_1_in_valid = PENetwork_11_io_to_pes_1_in_valid; // @[pe.scala 262:34]
  assign PE_1_io_data_1_in_bits = PENetwork_11_io_to_pes_1_in_bits; // @[pe.scala 262:34]
  assign PE_1_io_data_0_in_valid = PENetwork_1_io_to_pes_0_in_valid; // @[pe.scala 262:34]
  assign PE_1_io_data_0_in_bits = PENetwork_1_io_to_pes_0_in_bits; // @[pe.scala 262:34]
  assign PE_2_clock = clock;
  assign PE_2_reset = reset;
  assign PE_2_io_data_2_in_valid = PENetwork_26_io_to_pes_2_in_valid; // @[pe.scala 262:34]
  assign PE_2_io_data_2_in_bits = PENetwork_26_io_to_pes_2_in_bits; // @[pe.scala 262:34]
  assign PE_2_io_data_2_sig_stat2trans = PENetwork_26_io_to_pes_2_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_2_io_data_2_out_ready = PENetwork_26_io_to_pes_2_out_ready; // @[pe.scala 268:49]
  assign PE_2_io_data_1_in_valid = PENetwork_11_io_to_pes_2_in_valid; // @[pe.scala 262:34]
  assign PE_2_io_data_1_in_bits = PENetwork_11_io_to_pes_2_in_bits; // @[pe.scala 262:34]
  assign PE_2_io_data_0_in_valid = PENetwork_2_io_to_pes_0_in_valid; // @[pe.scala 262:34]
  assign PE_2_io_data_0_in_bits = PENetwork_2_io_to_pes_0_in_bits; // @[pe.scala 262:34]
  assign PE_3_clock = clock;
  assign PE_3_reset = reset;
  assign PE_3_io_data_2_in_valid = PENetwork_26_io_to_pes_3_in_valid; // @[pe.scala 262:34]
  assign PE_3_io_data_2_in_bits = PENetwork_26_io_to_pes_3_in_bits; // @[pe.scala 262:34]
  assign PE_3_io_data_2_sig_stat2trans = PENetwork_26_io_to_pes_3_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_3_io_data_2_out_ready = PENetwork_26_io_to_pes_3_out_ready; // @[pe.scala 268:49]
  assign PE_3_io_data_1_in_valid = PENetwork_11_io_to_pes_3_in_valid; // @[pe.scala 262:34]
  assign PE_3_io_data_1_in_bits = PENetwork_11_io_to_pes_3_in_bits; // @[pe.scala 262:34]
  assign PE_3_io_data_0_in_valid = PENetwork_3_io_to_pes_0_in_valid; // @[pe.scala 262:34]
  assign PE_3_io_data_0_in_bits = PENetwork_3_io_to_pes_0_in_bits; // @[pe.scala 262:34]
  assign PE_4_clock = clock;
  assign PE_4_reset = reset;
  assign PE_4_io_data_2_in_valid = PENetwork_26_io_to_pes_4_in_valid; // @[pe.scala 262:34]
  assign PE_4_io_data_2_in_bits = PENetwork_26_io_to_pes_4_in_bits; // @[pe.scala 262:34]
  assign PE_4_io_data_2_sig_stat2trans = PENetwork_26_io_to_pes_4_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_4_io_data_2_out_ready = PENetwork_26_io_to_pes_4_out_ready; // @[pe.scala 268:49]
  assign PE_4_io_data_1_in_valid = PENetwork_11_io_to_pes_4_in_valid; // @[pe.scala 262:34]
  assign PE_4_io_data_1_in_bits = PENetwork_11_io_to_pes_4_in_bits; // @[pe.scala 262:34]
  assign PE_4_io_data_0_in_valid = PENetwork_4_io_to_pes_0_in_valid; // @[pe.scala 262:34]
  assign PE_4_io_data_0_in_bits = PENetwork_4_io_to_pes_0_in_bits; // @[pe.scala 262:34]
  assign PE_5_clock = clock;
  assign PE_5_reset = reset;
  assign PE_5_io_data_2_in_valid = PENetwork_26_io_to_pes_5_in_valid; // @[pe.scala 262:34]
  assign PE_5_io_data_2_in_bits = PENetwork_26_io_to_pes_5_in_bits; // @[pe.scala 262:34]
  assign PE_5_io_data_2_sig_stat2trans = PENetwork_26_io_to_pes_5_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_5_io_data_2_out_ready = PENetwork_26_io_to_pes_5_out_ready; // @[pe.scala 268:49]
  assign PE_5_io_data_1_in_valid = PENetwork_11_io_to_pes_5_in_valid; // @[pe.scala 262:34]
  assign PE_5_io_data_1_in_bits = PENetwork_11_io_to_pes_5_in_bits; // @[pe.scala 262:34]
  assign PE_5_io_data_0_in_valid = PENetwork_5_io_to_pes_0_in_valid; // @[pe.scala 262:34]
  assign PE_5_io_data_0_in_bits = PENetwork_5_io_to_pes_0_in_bits; // @[pe.scala 262:34]
  assign PE_6_clock = clock;
  assign PE_6_reset = reset;
  assign PE_6_io_data_2_in_valid = PENetwork_26_io_to_pes_6_in_valid; // @[pe.scala 262:34]
  assign PE_6_io_data_2_in_bits = PENetwork_26_io_to_pes_6_in_bits; // @[pe.scala 262:34]
  assign PE_6_io_data_2_sig_stat2trans = PENetwork_26_io_to_pes_6_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_6_io_data_2_out_ready = PENetwork_26_io_to_pes_6_out_ready; // @[pe.scala 268:49]
  assign PE_6_io_data_1_in_valid = PENetwork_11_io_to_pes_6_in_valid; // @[pe.scala 262:34]
  assign PE_6_io_data_1_in_bits = PENetwork_11_io_to_pes_6_in_bits; // @[pe.scala 262:34]
  assign PE_6_io_data_0_in_valid = PENetwork_6_io_to_pes_0_in_valid; // @[pe.scala 262:34]
  assign PE_6_io_data_0_in_bits = PENetwork_6_io_to_pes_0_in_bits; // @[pe.scala 262:34]
  assign PE_7_clock = clock;
  assign PE_7_reset = reset;
  assign PE_7_io_data_2_in_valid = PENetwork_26_io_to_pes_7_in_valid; // @[pe.scala 262:34]
  assign PE_7_io_data_2_in_bits = PENetwork_26_io_to_pes_7_in_bits; // @[pe.scala 262:34]
  assign PE_7_io_data_2_sig_stat2trans = PENetwork_26_io_to_pes_7_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_7_io_data_2_out_ready = PENetwork_26_io_to_pes_7_out_ready; // @[pe.scala 268:49]
  assign PE_7_io_data_1_in_valid = PENetwork_11_io_to_pes_7_in_valid; // @[pe.scala 262:34]
  assign PE_7_io_data_1_in_bits = PENetwork_11_io_to_pes_7_in_bits; // @[pe.scala 262:34]
  assign PE_7_io_data_0_in_valid = PENetwork_7_io_to_pes_0_in_valid; // @[pe.scala 262:34]
  assign PE_7_io_data_0_in_bits = PENetwork_7_io_to_pes_0_in_bits; // @[pe.scala 262:34]
  assign PE_8_clock = clock;
  assign PE_8_reset = reset;
  assign PE_8_io_data_2_in_valid = PENetwork_26_io_to_pes_8_in_valid; // @[pe.scala 262:34]
  assign PE_8_io_data_2_in_bits = PENetwork_26_io_to_pes_8_in_bits; // @[pe.scala 262:34]
  assign PE_8_io_data_2_sig_stat2trans = PENetwork_26_io_to_pes_8_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_8_io_data_2_out_ready = PENetwork_26_io_to_pes_8_out_ready; // @[pe.scala 268:49]
  assign PE_8_io_data_1_in_valid = PENetwork_11_io_to_pes_8_in_valid; // @[pe.scala 262:34]
  assign PE_8_io_data_1_in_bits = PENetwork_11_io_to_pes_8_in_bits; // @[pe.scala 262:34]
  assign PE_8_io_data_0_in_valid = PENetwork_8_io_to_pes_0_in_valid; // @[pe.scala 262:34]
  assign PE_8_io_data_0_in_bits = PENetwork_8_io_to_pes_0_in_bits; // @[pe.scala 262:34]
  assign PE_9_clock = clock;
  assign PE_9_reset = reset;
  assign PE_9_io_data_2_in_valid = PENetwork_26_io_to_pes_9_in_valid; // @[pe.scala 262:34]
  assign PE_9_io_data_2_in_bits = PENetwork_26_io_to_pes_9_in_bits; // @[pe.scala 262:34]
  assign PE_9_io_data_2_sig_stat2trans = PENetwork_26_io_to_pes_9_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_9_io_data_2_out_ready = PENetwork_26_io_to_pes_9_out_ready; // @[pe.scala 268:49]
  assign PE_9_io_data_1_in_valid = PENetwork_11_io_to_pes_9_in_valid; // @[pe.scala 262:34]
  assign PE_9_io_data_1_in_bits = PENetwork_11_io_to_pes_9_in_bits; // @[pe.scala 262:34]
  assign PE_9_io_data_0_in_valid = PENetwork_9_io_to_pes_0_in_valid; // @[pe.scala 262:34]
  assign PE_9_io_data_0_in_bits = PENetwork_9_io_to_pes_0_in_bits; // @[pe.scala 262:34]
  assign PE_10_clock = clock;
  assign PE_10_reset = reset;
  assign PE_10_io_data_2_in_valid = PENetwork_26_io_to_pes_10_in_valid; // @[pe.scala 262:34]
  assign PE_10_io_data_2_in_bits = PENetwork_26_io_to_pes_10_in_bits; // @[pe.scala 262:34]
  assign PE_10_io_data_2_sig_stat2trans = PENetwork_26_io_to_pes_10_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_10_io_data_2_out_ready = 1'h1; // @[pe.scala 268:49]
  assign PE_10_io_data_1_in_valid = PENetwork_11_io_to_pes_10_in_valid; // @[pe.scala 262:34]
  assign PE_10_io_data_1_in_bits = PENetwork_11_io_to_pes_10_in_bits; // @[pe.scala 262:34]
  assign PE_10_io_data_0_in_valid = PENetwork_10_io_to_pes_0_in_valid; // @[pe.scala 262:34]
  assign PE_10_io_data_0_in_bits = PENetwork_10_io_to_pes_0_in_bits; // @[pe.scala 262:34]
  assign PE_11_clock = clock;
  assign PE_11_reset = reset;
  assign PE_11_io_data_2_in_valid = 1'h0; // @[pe.scala 262:34]
  assign PE_11_io_data_2_in_bits = 256'h0; // @[pe.scala 262:34]
  assign PE_11_io_data_2_sig_stat2trans = PENetwork_27_io_to_pes_0_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_11_io_data_2_out_ready = PENetwork_27_io_to_pes_0_out_ready; // @[pe.scala 268:49]
  assign PE_11_io_data_1_in_valid = PENetwork_12_io_to_pes_0_in_valid; // @[pe.scala 262:34]
  assign PE_11_io_data_1_in_bits = PENetwork_12_io_to_pes_0_in_bits; // @[pe.scala 262:34]
  assign PE_11_io_data_0_in_valid = PENetwork_io_to_pes_1_in_valid; // @[pe.scala 262:34]
  assign PE_11_io_data_0_in_bits = PENetwork_io_to_pes_1_in_bits; // @[pe.scala 262:34]
  assign PE_12_clock = clock;
  assign PE_12_reset = reset;
  assign PE_12_io_data_2_in_valid = PENetwork_27_io_to_pes_1_in_valid; // @[pe.scala 262:34]
  assign PE_12_io_data_2_in_bits = PENetwork_27_io_to_pes_1_in_bits; // @[pe.scala 262:34]
  assign PE_12_io_data_2_sig_stat2trans = PENetwork_27_io_to_pes_1_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_12_io_data_2_out_ready = PENetwork_27_io_to_pes_1_out_ready; // @[pe.scala 268:49]
  assign PE_12_io_data_1_in_valid = PENetwork_12_io_to_pes_1_in_valid; // @[pe.scala 262:34]
  assign PE_12_io_data_1_in_bits = PENetwork_12_io_to_pes_1_in_bits; // @[pe.scala 262:34]
  assign PE_12_io_data_0_in_valid = PENetwork_1_io_to_pes_1_in_valid; // @[pe.scala 262:34]
  assign PE_12_io_data_0_in_bits = PENetwork_1_io_to_pes_1_in_bits; // @[pe.scala 262:34]
  assign PE_13_clock = clock;
  assign PE_13_reset = reset;
  assign PE_13_io_data_2_in_valid = PENetwork_27_io_to_pes_2_in_valid; // @[pe.scala 262:34]
  assign PE_13_io_data_2_in_bits = PENetwork_27_io_to_pes_2_in_bits; // @[pe.scala 262:34]
  assign PE_13_io_data_2_sig_stat2trans = PENetwork_27_io_to_pes_2_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_13_io_data_2_out_ready = PENetwork_27_io_to_pes_2_out_ready; // @[pe.scala 268:49]
  assign PE_13_io_data_1_in_valid = PENetwork_12_io_to_pes_2_in_valid; // @[pe.scala 262:34]
  assign PE_13_io_data_1_in_bits = PENetwork_12_io_to_pes_2_in_bits; // @[pe.scala 262:34]
  assign PE_13_io_data_0_in_valid = PENetwork_2_io_to_pes_1_in_valid; // @[pe.scala 262:34]
  assign PE_13_io_data_0_in_bits = PENetwork_2_io_to_pes_1_in_bits; // @[pe.scala 262:34]
  assign PE_14_clock = clock;
  assign PE_14_reset = reset;
  assign PE_14_io_data_2_in_valid = PENetwork_27_io_to_pes_3_in_valid; // @[pe.scala 262:34]
  assign PE_14_io_data_2_in_bits = PENetwork_27_io_to_pes_3_in_bits; // @[pe.scala 262:34]
  assign PE_14_io_data_2_sig_stat2trans = PENetwork_27_io_to_pes_3_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_14_io_data_2_out_ready = PENetwork_27_io_to_pes_3_out_ready; // @[pe.scala 268:49]
  assign PE_14_io_data_1_in_valid = PENetwork_12_io_to_pes_3_in_valid; // @[pe.scala 262:34]
  assign PE_14_io_data_1_in_bits = PENetwork_12_io_to_pes_3_in_bits; // @[pe.scala 262:34]
  assign PE_14_io_data_0_in_valid = PENetwork_3_io_to_pes_1_in_valid; // @[pe.scala 262:34]
  assign PE_14_io_data_0_in_bits = PENetwork_3_io_to_pes_1_in_bits; // @[pe.scala 262:34]
  assign PE_15_clock = clock;
  assign PE_15_reset = reset;
  assign PE_15_io_data_2_in_valid = PENetwork_27_io_to_pes_4_in_valid; // @[pe.scala 262:34]
  assign PE_15_io_data_2_in_bits = PENetwork_27_io_to_pes_4_in_bits; // @[pe.scala 262:34]
  assign PE_15_io_data_2_sig_stat2trans = PENetwork_27_io_to_pes_4_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_15_io_data_2_out_ready = PENetwork_27_io_to_pes_4_out_ready; // @[pe.scala 268:49]
  assign PE_15_io_data_1_in_valid = PENetwork_12_io_to_pes_4_in_valid; // @[pe.scala 262:34]
  assign PE_15_io_data_1_in_bits = PENetwork_12_io_to_pes_4_in_bits; // @[pe.scala 262:34]
  assign PE_15_io_data_0_in_valid = PENetwork_4_io_to_pes_1_in_valid; // @[pe.scala 262:34]
  assign PE_15_io_data_0_in_bits = PENetwork_4_io_to_pes_1_in_bits; // @[pe.scala 262:34]
  assign PE_16_clock = clock;
  assign PE_16_reset = reset;
  assign PE_16_io_data_2_in_valid = PENetwork_27_io_to_pes_5_in_valid; // @[pe.scala 262:34]
  assign PE_16_io_data_2_in_bits = PENetwork_27_io_to_pes_5_in_bits; // @[pe.scala 262:34]
  assign PE_16_io_data_2_sig_stat2trans = PENetwork_27_io_to_pes_5_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_16_io_data_2_out_ready = PENetwork_27_io_to_pes_5_out_ready; // @[pe.scala 268:49]
  assign PE_16_io_data_1_in_valid = PENetwork_12_io_to_pes_5_in_valid; // @[pe.scala 262:34]
  assign PE_16_io_data_1_in_bits = PENetwork_12_io_to_pes_5_in_bits; // @[pe.scala 262:34]
  assign PE_16_io_data_0_in_valid = PENetwork_5_io_to_pes_1_in_valid; // @[pe.scala 262:34]
  assign PE_16_io_data_0_in_bits = PENetwork_5_io_to_pes_1_in_bits; // @[pe.scala 262:34]
  assign PE_17_clock = clock;
  assign PE_17_reset = reset;
  assign PE_17_io_data_2_in_valid = PENetwork_27_io_to_pes_6_in_valid; // @[pe.scala 262:34]
  assign PE_17_io_data_2_in_bits = PENetwork_27_io_to_pes_6_in_bits; // @[pe.scala 262:34]
  assign PE_17_io_data_2_sig_stat2trans = PENetwork_27_io_to_pes_6_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_17_io_data_2_out_ready = PENetwork_27_io_to_pes_6_out_ready; // @[pe.scala 268:49]
  assign PE_17_io_data_1_in_valid = PENetwork_12_io_to_pes_6_in_valid; // @[pe.scala 262:34]
  assign PE_17_io_data_1_in_bits = PENetwork_12_io_to_pes_6_in_bits; // @[pe.scala 262:34]
  assign PE_17_io_data_0_in_valid = PENetwork_6_io_to_pes_1_in_valid; // @[pe.scala 262:34]
  assign PE_17_io_data_0_in_bits = PENetwork_6_io_to_pes_1_in_bits; // @[pe.scala 262:34]
  assign PE_18_clock = clock;
  assign PE_18_reset = reset;
  assign PE_18_io_data_2_in_valid = PENetwork_27_io_to_pes_7_in_valid; // @[pe.scala 262:34]
  assign PE_18_io_data_2_in_bits = PENetwork_27_io_to_pes_7_in_bits; // @[pe.scala 262:34]
  assign PE_18_io_data_2_sig_stat2trans = PENetwork_27_io_to_pes_7_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_18_io_data_2_out_ready = PENetwork_27_io_to_pes_7_out_ready; // @[pe.scala 268:49]
  assign PE_18_io_data_1_in_valid = PENetwork_12_io_to_pes_7_in_valid; // @[pe.scala 262:34]
  assign PE_18_io_data_1_in_bits = PENetwork_12_io_to_pes_7_in_bits; // @[pe.scala 262:34]
  assign PE_18_io_data_0_in_valid = PENetwork_7_io_to_pes_1_in_valid; // @[pe.scala 262:34]
  assign PE_18_io_data_0_in_bits = PENetwork_7_io_to_pes_1_in_bits; // @[pe.scala 262:34]
  assign PE_19_clock = clock;
  assign PE_19_reset = reset;
  assign PE_19_io_data_2_in_valid = PENetwork_27_io_to_pes_8_in_valid; // @[pe.scala 262:34]
  assign PE_19_io_data_2_in_bits = PENetwork_27_io_to_pes_8_in_bits; // @[pe.scala 262:34]
  assign PE_19_io_data_2_sig_stat2trans = PENetwork_27_io_to_pes_8_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_19_io_data_2_out_ready = PENetwork_27_io_to_pes_8_out_ready; // @[pe.scala 268:49]
  assign PE_19_io_data_1_in_valid = PENetwork_12_io_to_pes_8_in_valid; // @[pe.scala 262:34]
  assign PE_19_io_data_1_in_bits = PENetwork_12_io_to_pes_8_in_bits; // @[pe.scala 262:34]
  assign PE_19_io_data_0_in_valid = PENetwork_8_io_to_pes_1_in_valid; // @[pe.scala 262:34]
  assign PE_19_io_data_0_in_bits = PENetwork_8_io_to_pes_1_in_bits; // @[pe.scala 262:34]
  assign PE_20_clock = clock;
  assign PE_20_reset = reset;
  assign PE_20_io_data_2_in_valid = PENetwork_27_io_to_pes_9_in_valid; // @[pe.scala 262:34]
  assign PE_20_io_data_2_in_bits = PENetwork_27_io_to_pes_9_in_bits; // @[pe.scala 262:34]
  assign PE_20_io_data_2_sig_stat2trans = PENetwork_27_io_to_pes_9_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_20_io_data_2_out_ready = PENetwork_27_io_to_pes_9_out_ready; // @[pe.scala 268:49]
  assign PE_20_io_data_1_in_valid = PENetwork_12_io_to_pes_9_in_valid; // @[pe.scala 262:34]
  assign PE_20_io_data_1_in_bits = PENetwork_12_io_to_pes_9_in_bits; // @[pe.scala 262:34]
  assign PE_20_io_data_0_in_valid = PENetwork_9_io_to_pes_1_in_valid; // @[pe.scala 262:34]
  assign PE_20_io_data_0_in_bits = PENetwork_9_io_to_pes_1_in_bits; // @[pe.scala 262:34]
  assign PE_21_clock = clock;
  assign PE_21_reset = reset;
  assign PE_21_io_data_2_in_valid = PENetwork_27_io_to_pes_10_in_valid; // @[pe.scala 262:34]
  assign PE_21_io_data_2_in_bits = PENetwork_27_io_to_pes_10_in_bits; // @[pe.scala 262:34]
  assign PE_21_io_data_2_sig_stat2trans = PENetwork_27_io_to_pes_10_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_21_io_data_2_out_ready = 1'h1; // @[pe.scala 268:49]
  assign PE_21_io_data_1_in_valid = PENetwork_12_io_to_pes_10_in_valid; // @[pe.scala 262:34]
  assign PE_21_io_data_1_in_bits = PENetwork_12_io_to_pes_10_in_bits; // @[pe.scala 262:34]
  assign PE_21_io_data_0_in_valid = PENetwork_10_io_to_pes_1_in_valid; // @[pe.scala 262:34]
  assign PE_21_io_data_0_in_bits = PENetwork_10_io_to_pes_1_in_bits; // @[pe.scala 262:34]
  assign PE_22_clock = clock;
  assign PE_22_reset = reset;
  assign PE_22_io_data_2_in_valid = 1'h0; // @[pe.scala 262:34]
  assign PE_22_io_data_2_in_bits = 256'h0; // @[pe.scala 262:34]
  assign PE_22_io_data_2_sig_stat2trans = PENetwork_28_io_to_pes_0_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_22_io_data_2_out_ready = PENetwork_28_io_to_pes_0_out_ready; // @[pe.scala 268:49]
  assign PE_22_io_data_1_in_valid = PENetwork_13_io_to_pes_0_in_valid; // @[pe.scala 262:34]
  assign PE_22_io_data_1_in_bits = PENetwork_13_io_to_pes_0_in_bits; // @[pe.scala 262:34]
  assign PE_22_io_data_0_in_valid = PENetwork_io_to_pes_2_in_valid; // @[pe.scala 262:34]
  assign PE_22_io_data_0_in_bits = PENetwork_io_to_pes_2_in_bits; // @[pe.scala 262:34]
  assign PE_23_clock = clock;
  assign PE_23_reset = reset;
  assign PE_23_io_data_2_in_valid = PENetwork_28_io_to_pes_1_in_valid; // @[pe.scala 262:34]
  assign PE_23_io_data_2_in_bits = PENetwork_28_io_to_pes_1_in_bits; // @[pe.scala 262:34]
  assign PE_23_io_data_2_sig_stat2trans = PENetwork_28_io_to_pes_1_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_23_io_data_2_out_ready = PENetwork_28_io_to_pes_1_out_ready; // @[pe.scala 268:49]
  assign PE_23_io_data_1_in_valid = PENetwork_13_io_to_pes_1_in_valid; // @[pe.scala 262:34]
  assign PE_23_io_data_1_in_bits = PENetwork_13_io_to_pes_1_in_bits; // @[pe.scala 262:34]
  assign PE_23_io_data_0_in_valid = PENetwork_1_io_to_pes_2_in_valid; // @[pe.scala 262:34]
  assign PE_23_io_data_0_in_bits = PENetwork_1_io_to_pes_2_in_bits; // @[pe.scala 262:34]
  assign PE_24_clock = clock;
  assign PE_24_reset = reset;
  assign PE_24_io_data_2_in_valid = PENetwork_28_io_to_pes_2_in_valid; // @[pe.scala 262:34]
  assign PE_24_io_data_2_in_bits = PENetwork_28_io_to_pes_2_in_bits; // @[pe.scala 262:34]
  assign PE_24_io_data_2_sig_stat2trans = PENetwork_28_io_to_pes_2_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_24_io_data_2_out_ready = PENetwork_28_io_to_pes_2_out_ready; // @[pe.scala 268:49]
  assign PE_24_io_data_1_in_valid = PENetwork_13_io_to_pes_2_in_valid; // @[pe.scala 262:34]
  assign PE_24_io_data_1_in_bits = PENetwork_13_io_to_pes_2_in_bits; // @[pe.scala 262:34]
  assign PE_24_io_data_0_in_valid = PENetwork_2_io_to_pes_2_in_valid; // @[pe.scala 262:34]
  assign PE_24_io_data_0_in_bits = PENetwork_2_io_to_pes_2_in_bits; // @[pe.scala 262:34]
  assign PE_25_clock = clock;
  assign PE_25_reset = reset;
  assign PE_25_io_data_2_in_valid = PENetwork_28_io_to_pes_3_in_valid; // @[pe.scala 262:34]
  assign PE_25_io_data_2_in_bits = PENetwork_28_io_to_pes_3_in_bits; // @[pe.scala 262:34]
  assign PE_25_io_data_2_sig_stat2trans = PENetwork_28_io_to_pes_3_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_25_io_data_2_out_ready = PENetwork_28_io_to_pes_3_out_ready; // @[pe.scala 268:49]
  assign PE_25_io_data_1_in_valid = PENetwork_13_io_to_pes_3_in_valid; // @[pe.scala 262:34]
  assign PE_25_io_data_1_in_bits = PENetwork_13_io_to_pes_3_in_bits; // @[pe.scala 262:34]
  assign PE_25_io_data_0_in_valid = PENetwork_3_io_to_pes_2_in_valid; // @[pe.scala 262:34]
  assign PE_25_io_data_0_in_bits = PENetwork_3_io_to_pes_2_in_bits; // @[pe.scala 262:34]
  assign PE_26_clock = clock;
  assign PE_26_reset = reset;
  assign PE_26_io_data_2_in_valid = PENetwork_28_io_to_pes_4_in_valid; // @[pe.scala 262:34]
  assign PE_26_io_data_2_in_bits = PENetwork_28_io_to_pes_4_in_bits; // @[pe.scala 262:34]
  assign PE_26_io_data_2_sig_stat2trans = PENetwork_28_io_to_pes_4_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_26_io_data_2_out_ready = PENetwork_28_io_to_pes_4_out_ready; // @[pe.scala 268:49]
  assign PE_26_io_data_1_in_valid = PENetwork_13_io_to_pes_4_in_valid; // @[pe.scala 262:34]
  assign PE_26_io_data_1_in_bits = PENetwork_13_io_to_pes_4_in_bits; // @[pe.scala 262:34]
  assign PE_26_io_data_0_in_valid = PENetwork_4_io_to_pes_2_in_valid; // @[pe.scala 262:34]
  assign PE_26_io_data_0_in_bits = PENetwork_4_io_to_pes_2_in_bits; // @[pe.scala 262:34]
  assign PE_27_clock = clock;
  assign PE_27_reset = reset;
  assign PE_27_io_data_2_in_valid = PENetwork_28_io_to_pes_5_in_valid; // @[pe.scala 262:34]
  assign PE_27_io_data_2_in_bits = PENetwork_28_io_to_pes_5_in_bits; // @[pe.scala 262:34]
  assign PE_27_io_data_2_sig_stat2trans = PENetwork_28_io_to_pes_5_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_27_io_data_2_out_ready = PENetwork_28_io_to_pes_5_out_ready; // @[pe.scala 268:49]
  assign PE_27_io_data_1_in_valid = PENetwork_13_io_to_pes_5_in_valid; // @[pe.scala 262:34]
  assign PE_27_io_data_1_in_bits = PENetwork_13_io_to_pes_5_in_bits; // @[pe.scala 262:34]
  assign PE_27_io_data_0_in_valid = PENetwork_5_io_to_pes_2_in_valid; // @[pe.scala 262:34]
  assign PE_27_io_data_0_in_bits = PENetwork_5_io_to_pes_2_in_bits; // @[pe.scala 262:34]
  assign PE_28_clock = clock;
  assign PE_28_reset = reset;
  assign PE_28_io_data_2_in_valid = PENetwork_28_io_to_pes_6_in_valid; // @[pe.scala 262:34]
  assign PE_28_io_data_2_in_bits = PENetwork_28_io_to_pes_6_in_bits; // @[pe.scala 262:34]
  assign PE_28_io_data_2_sig_stat2trans = PENetwork_28_io_to_pes_6_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_28_io_data_2_out_ready = PENetwork_28_io_to_pes_6_out_ready; // @[pe.scala 268:49]
  assign PE_28_io_data_1_in_valid = PENetwork_13_io_to_pes_6_in_valid; // @[pe.scala 262:34]
  assign PE_28_io_data_1_in_bits = PENetwork_13_io_to_pes_6_in_bits; // @[pe.scala 262:34]
  assign PE_28_io_data_0_in_valid = PENetwork_6_io_to_pes_2_in_valid; // @[pe.scala 262:34]
  assign PE_28_io_data_0_in_bits = PENetwork_6_io_to_pes_2_in_bits; // @[pe.scala 262:34]
  assign PE_29_clock = clock;
  assign PE_29_reset = reset;
  assign PE_29_io_data_2_in_valid = PENetwork_28_io_to_pes_7_in_valid; // @[pe.scala 262:34]
  assign PE_29_io_data_2_in_bits = PENetwork_28_io_to_pes_7_in_bits; // @[pe.scala 262:34]
  assign PE_29_io_data_2_sig_stat2trans = PENetwork_28_io_to_pes_7_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_29_io_data_2_out_ready = PENetwork_28_io_to_pes_7_out_ready; // @[pe.scala 268:49]
  assign PE_29_io_data_1_in_valid = PENetwork_13_io_to_pes_7_in_valid; // @[pe.scala 262:34]
  assign PE_29_io_data_1_in_bits = PENetwork_13_io_to_pes_7_in_bits; // @[pe.scala 262:34]
  assign PE_29_io_data_0_in_valid = PENetwork_7_io_to_pes_2_in_valid; // @[pe.scala 262:34]
  assign PE_29_io_data_0_in_bits = PENetwork_7_io_to_pes_2_in_bits; // @[pe.scala 262:34]
  assign PE_30_clock = clock;
  assign PE_30_reset = reset;
  assign PE_30_io_data_2_in_valid = PENetwork_28_io_to_pes_8_in_valid; // @[pe.scala 262:34]
  assign PE_30_io_data_2_in_bits = PENetwork_28_io_to_pes_8_in_bits; // @[pe.scala 262:34]
  assign PE_30_io_data_2_sig_stat2trans = PENetwork_28_io_to_pes_8_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_30_io_data_2_out_ready = PENetwork_28_io_to_pes_8_out_ready; // @[pe.scala 268:49]
  assign PE_30_io_data_1_in_valid = PENetwork_13_io_to_pes_8_in_valid; // @[pe.scala 262:34]
  assign PE_30_io_data_1_in_bits = PENetwork_13_io_to_pes_8_in_bits; // @[pe.scala 262:34]
  assign PE_30_io_data_0_in_valid = PENetwork_8_io_to_pes_2_in_valid; // @[pe.scala 262:34]
  assign PE_30_io_data_0_in_bits = PENetwork_8_io_to_pes_2_in_bits; // @[pe.scala 262:34]
  assign PE_31_clock = clock;
  assign PE_31_reset = reset;
  assign PE_31_io_data_2_in_valid = PENetwork_28_io_to_pes_9_in_valid; // @[pe.scala 262:34]
  assign PE_31_io_data_2_in_bits = PENetwork_28_io_to_pes_9_in_bits; // @[pe.scala 262:34]
  assign PE_31_io_data_2_sig_stat2trans = PENetwork_28_io_to_pes_9_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_31_io_data_2_out_ready = PENetwork_28_io_to_pes_9_out_ready; // @[pe.scala 268:49]
  assign PE_31_io_data_1_in_valid = PENetwork_13_io_to_pes_9_in_valid; // @[pe.scala 262:34]
  assign PE_31_io_data_1_in_bits = PENetwork_13_io_to_pes_9_in_bits; // @[pe.scala 262:34]
  assign PE_31_io_data_0_in_valid = PENetwork_9_io_to_pes_2_in_valid; // @[pe.scala 262:34]
  assign PE_31_io_data_0_in_bits = PENetwork_9_io_to_pes_2_in_bits; // @[pe.scala 262:34]
  assign PE_32_clock = clock;
  assign PE_32_reset = reset;
  assign PE_32_io_data_2_in_valid = PENetwork_28_io_to_pes_10_in_valid; // @[pe.scala 262:34]
  assign PE_32_io_data_2_in_bits = PENetwork_28_io_to_pes_10_in_bits; // @[pe.scala 262:34]
  assign PE_32_io_data_2_sig_stat2trans = PENetwork_28_io_to_pes_10_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_32_io_data_2_out_ready = 1'h1; // @[pe.scala 268:49]
  assign PE_32_io_data_1_in_valid = PENetwork_13_io_to_pes_10_in_valid; // @[pe.scala 262:34]
  assign PE_32_io_data_1_in_bits = PENetwork_13_io_to_pes_10_in_bits; // @[pe.scala 262:34]
  assign PE_32_io_data_0_in_valid = PENetwork_10_io_to_pes_2_in_valid; // @[pe.scala 262:34]
  assign PE_32_io_data_0_in_bits = PENetwork_10_io_to_pes_2_in_bits; // @[pe.scala 262:34]
  assign PE_33_clock = clock;
  assign PE_33_reset = reset;
  assign PE_33_io_data_2_in_valid = 1'h0; // @[pe.scala 262:34]
  assign PE_33_io_data_2_in_bits = 256'h0; // @[pe.scala 262:34]
  assign PE_33_io_data_2_sig_stat2trans = PENetwork_29_io_to_pes_0_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_33_io_data_2_out_ready = PENetwork_29_io_to_pes_0_out_ready; // @[pe.scala 268:49]
  assign PE_33_io_data_1_in_valid = PENetwork_14_io_to_pes_0_in_valid; // @[pe.scala 262:34]
  assign PE_33_io_data_1_in_bits = PENetwork_14_io_to_pes_0_in_bits; // @[pe.scala 262:34]
  assign PE_33_io_data_0_in_valid = PENetwork_io_to_pes_3_in_valid; // @[pe.scala 262:34]
  assign PE_33_io_data_0_in_bits = PENetwork_io_to_pes_3_in_bits; // @[pe.scala 262:34]
  assign PE_34_clock = clock;
  assign PE_34_reset = reset;
  assign PE_34_io_data_2_in_valid = PENetwork_29_io_to_pes_1_in_valid; // @[pe.scala 262:34]
  assign PE_34_io_data_2_in_bits = PENetwork_29_io_to_pes_1_in_bits; // @[pe.scala 262:34]
  assign PE_34_io_data_2_sig_stat2trans = PENetwork_29_io_to_pes_1_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_34_io_data_2_out_ready = PENetwork_29_io_to_pes_1_out_ready; // @[pe.scala 268:49]
  assign PE_34_io_data_1_in_valid = PENetwork_14_io_to_pes_1_in_valid; // @[pe.scala 262:34]
  assign PE_34_io_data_1_in_bits = PENetwork_14_io_to_pes_1_in_bits; // @[pe.scala 262:34]
  assign PE_34_io_data_0_in_valid = PENetwork_1_io_to_pes_3_in_valid; // @[pe.scala 262:34]
  assign PE_34_io_data_0_in_bits = PENetwork_1_io_to_pes_3_in_bits; // @[pe.scala 262:34]
  assign PE_35_clock = clock;
  assign PE_35_reset = reset;
  assign PE_35_io_data_2_in_valid = PENetwork_29_io_to_pes_2_in_valid; // @[pe.scala 262:34]
  assign PE_35_io_data_2_in_bits = PENetwork_29_io_to_pes_2_in_bits; // @[pe.scala 262:34]
  assign PE_35_io_data_2_sig_stat2trans = PENetwork_29_io_to_pes_2_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_35_io_data_2_out_ready = PENetwork_29_io_to_pes_2_out_ready; // @[pe.scala 268:49]
  assign PE_35_io_data_1_in_valid = PENetwork_14_io_to_pes_2_in_valid; // @[pe.scala 262:34]
  assign PE_35_io_data_1_in_bits = PENetwork_14_io_to_pes_2_in_bits; // @[pe.scala 262:34]
  assign PE_35_io_data_0_in_valid = PENetwork_2_io_to_pes_3_in_valid; // @[pe.scala 262:34]
  assign PE_35_io_data_0_in_bits = PENetwork_2_io_to_pes_3_in_bits; // @[pe.scala 262:34]
  assign PE_36_clock = clock;
  assign PE_36_reset = reset;
  assign PE_36_io_data_2_in_valid = PENetwork_29_io_to_pes_3_in_valid; // @[pe.scala 262:34]
  assign PE_36_io_data_2_in_bits = PENetwork_29_io_to_pes_3_in_bits; // @[pe.scala 262:34]
  assign PE_36_io_data_2_sig_stat2trans = PENetwork_29_io_to_pes_3_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_36_io_data_2_out_ready = PENetwork_29_io_to_pes_3_out_ready; // @[pe.scala 268:49]
  assign PE_36_io_data_1_in_valid = PENetwork_14_io_to_pes_3_in_valid; // @[pe.scala 262:34]
  assign PE_36_io_data_1_in_bits = PENetwork_14_io_to_pes_3_in_bits; // @[pe.scala 262:34]
  assign PE_36_io_data_0_in_valid = PENetwork_3_io_to_pes_3_in_valid; // @[pe.scala 262:34]
  assign PE_36_io_data_0_in_bits = PENetwork_3_io_to_pes_3_in_bits; // @[pe.scala 262:34]
  assign PE_37_clock = clock;
  assign PE_37_reset = reset;
  assign PE_37_io_data_2_in_valid = PENetwork_29_io_to_pes_4_in_valid; // @[pe.scala 262:34]
  assign PE_37_io_data_2_in_bits = PENetwork_29_io_to_pes_4_in_bits; // @[pe.scala 262:34]
  assign PE_37_io_data_2_sig_stat2trans = PENetwork_29_io_to_pes_4_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_37_io_data_2_out_ready = PENetwork_29_io_to_pes_4_out_ready; // @[pe.scala 268:49]
  assign PE_37_io_data_1_in_valid = PENetwork_14_io_to_pes_4_in_valid; // @[pe.scala 262:34]
  assign PE_37_io_data_1_in_bits = PENetwork_14_io_to_pes_4_in_bits; // @[pe.scala 262:34]
  assign PE_37_io_data_0_in_valid = PENetwork_4_io_to_pes_3_in_valid; // @[pe.scala 262:34]
  assign PE_37_io_data_0_in_bits = PENetwork_4_io_to_pes_3_in_bits; // @[pe.scala 262:34]
  assign PE_38_clock = clock;
  assign PE_38_reset = reset;
  assign PE_38_io_data_2_in_valid = PENetwork_29_io_to_pes_5_in_valid; // @[pe.scala 262:34]
  assign PE_38_io_data_2_in_bits = PENetwork_29_io_to_pes_5_in_bits; // @[pe.scala 262:34]
  assign PE_38_io_data_2_sig_stat2trans = PENetwork_29_io_to_pes_5_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_38_io_data_2_out_ready = PENetwork_29_io_to_pes_5_out_ready; // @[pe.scala 268:49]
  assign PE_38_io_data_1_in_valid = PENetwork_14_io_to_pes_5_in_valid; // @[pe.scala 262:34]
  assign PE_38_io_data_1_in_bits = PENetwork_14_io_to_pes_5_in_bits; // @[pe.scala 262:34]
  assign PE_38_io_data_0_in_valid = PENetwork_5_io_to_pes_3_in_valid; // @[pe.scala 262:34]
  assign PE_38_io_data_0_in_bits = PENetwork_5_io_to_pes_3_in_bits; // @[pe.scala 262:34]
  assign PE_39_clock = clock;
  assign PE_39_reset = reset;
  assign PE_39_io_data_2_in_valid = PENetwork_29_io_to_pes_6_in_valid; // @[pe.scala 262:34]
  assign PE_39_io_data_2_in_bits = PENetwork_29_io_to_pes_6_in_bits; // @[pe.scala 262:34]
  assign PE_39_io_data_2_sig_stat2trans = PENetwork_29_io_to_pes_6_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_39_io_data_2_out_ready = PENetwork_29_io_to_pes_6_out_ready; // @[pe.scala 268:49]
  assign PE_39_io_data_1_in_valid = PENetwork_14_io_to_pes_6_in_valid; // @[pe.scala 262:34]
  assign PE_39_io_data_1_in_bits = PENetwork_14_io_to_pes_6_in_bits; // @[pe.scala 262:34]
  assign PE_39_io_data_0_in_valid = PENetwork_6_io_to_pes_3_in_valid; // @[pe.scala 262:34]
  assign PE_39_io_data_0_in_bits = PENetwork_6_io_to_pes_3_in_bits; // @[pe.scala 262:34]
  assign PE_40_clock = clock;
  assign PE_40_reset = reset;
  assign PE_40_io_data_2_in_valid = PENetwork_29_io_to_pes_7_in_valid; // @[pe.scala 262:34]
  assign PE_40_io_data_2_in_bits = PENetwork_29_io_to_pes_7_in_bits; // @[pe.scala 262:34]
  assign PE_40_io_data_2_sig_stat2trans = PENetwork_29_io_to_pes_7_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_40_io_data_2_out_ready = PENetwork_29_io_to_pes_7_out_ready; // @[pe.scala 268:49]
  assign PE_40_io_data_1_in_valid = PENetwork_14_io_to_pes_7_in_valid; // @[pe.scala 262:34]
  assign PE_40_io_data_1_in_bits = PENetwork_14_io_to_pes_7_in_bits; // @[pe.scala 262:34]
  assign PE_40_io_data_0_in_valid = PENetwork_7_io_to_pes_3_in_valid; // @[pe.scala 262:34]
  assign PE_40_io_data_0_in_bits = PENetwork_7_io_to_pes_3_in_bits; // @[pe.scala 262:34]
  assign PE_41_clock = clock;
  assign PE_41_reset = reset;
  assign PE_41_io_data_2_in_valid = PENetwork_29_io_to_pes_8_in_valid; // @[pe.scala 262:34]
  assign PE_41_io_data_2_in_bits = PENetwork_29_io_to_pes_8_in_bits; // @[pe.scala 262:34]
  assign PE_41_io_data_2_sig_stat2trans = PENetwork_29_io_to_pes_8_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_41_io_data_2_out_ready = PENetwork_29_io_to_pes_8_out_ready; // @[pe.scala 268:49]
  assign PE_41_io_data_1_in_valid = PENetwork_14_io_to_pes_8_in_valid; // @[pe.scala 262:34]
  assign PE_41_io_data_1_in_bits = PENetwork_14_io_to_pes_8_in_bits; // @[pe.scala 262:34]
  assign PE_41_io_data_0_in_valid = PENetwork_8_io_to_pes_3_in_valid; // @[pe.scala 262:34]
  assign PE_41_io_data_0_in_bits = PENetwork_8_io_to_pes_3_in_bits; // @[pe.scala 262:34]
  assign PE_42_clock = clock;
  assign PE_42_reset = reset;
  assign PE_42_io_data_2_in_valid = PENetwork_29_io_to_pes_9_in_valid; // @[pe.scala 262:34]
  assign PE_42_io_data_2_in_bits = PENetwork_29_io_to_pes_9_in_bits; // @[pe.scala 262:34]
  assign PE_42_io_data_2_sig_stat2trans = PENetwork_29_io_to_pes_9_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_42_io_data_2_out_ready = PENetwork_29_io_to_pes_9_out_ready; // @[pe.scala 268:49]
  assign PE_42_io_data_1_in_valid = PENetwork_14_io_to_pes_9_in_valid; // @[pe.scala 262:34]
  assign PE_42_io_data_1_in_bits = PENetwork_14_io_to_pes_9_in_bits; // @[pe.scala 262:34]
  assign PE_42_io_data_0_in_valid = PENetwork_9_io_to_pes_3_in_valid; // @[pe.scala 262:34]
  assign PE_42_io_data_0_in_bits = PENetwork_9_io_to_pes_3_in_bits; // @[pe.scala 262:34]
  assign PE_43_clock = clock;
  assign PE_43_reset = reset;
  assign PE_43_io_data_2_in_valid = PENetwork_29_io_to_pes_10_in_valid; // @[pe.scala 262:34]
  assign PE_43_io_data_2_in_bits = PENetwork_29_io_to_pes_10_in_bits; // @[pe.scala 262:34]
  assign PE_43_io_data_2_sig_stat2trans = PENetwork_29_io_to_pes_10_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_43_io_data_2_out_ready = 1'h1; // @[pe.scala 268:49]
  assign PE_43_io_data_1_in_valid = PENetwork_14_io_to_pes_10_in_valid; // @[pe.scala 262:34]
  assign PE_43_io_data_1_in_bits = PENetwork_14_io_to_pes_10_in_bits; // @[pe.scala 262:34]
  assign PE_43_io_data_0_in_valid = PENetwork_10_io_to_pes_3_in_valid; // @[pe.scala 262:34]
  assign PE_43_io_data_0_in_bits = PENetwork_10_io_to_pes_3_in_bits; // @[pe.scala 262:34]
  assign PE_44_clock = clock;
  assign PE_44_reset = reset;
  assign PE_44_io_data_2_in_valid = 1'h0; // @[pe.scala 262:34]
  assign PE_44_io_data_2_in_bits = 256'h0; // @[pe.scala 262:34]
  assign PE_44_io_data_2_sig_stat2trans = PENetwork_30_io_to_pes_0_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_44_io_data_2_out_ready = PENetwork_30_io_to_pes_0_out_ready; // @[pe.scala 268:49]
  assign PE_44_io_data_1_in_valid = PENetwork_15_io_to_pes_0_in_valid; // @[pe.scala 262:34]
  assign PE_44_io_data_1_in_bits = PENetwork_15_io_to_pes_0_in_bits; // @[pe.scala 262:34]
  assign PE_44_io_data_0_in_valid = PENetwork_io_to_pes_4_in_valid; // @[pe.scala 262:34]
  assign PE_44_io_data_0_in_bits = PENetwork_io_to_pes_4_in_bits; // @[pe.scala 262:34]
  assign PE_45_clock = clock;
  assign PE_45_reset = reset;
  assign PE_45_io_data_2_in_valid = PENetwork_30_io_to_pes_1_in_valid; // @[pe.scala 262:34]
  assign PE_45_io_data_2_in_bits = PENetwork_30_io_to_pes_1_in_bits; // @[pe.scala 262:34]
  assign PE_45_io_data_2_sig_stat2trans = PENetwork_30_io_to_pes_1_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_45_io_data_2_out_ready = PENetwork_30_io_to_pes_1_out_ready; // @[pe.scala 268:49]
  assign PE_45_io_data_1_in_valid = PENetwork_15_io_to_pes_1_in_valid; // @[pe.scala 262:34]
  assign PE_45_io_data_1_in_bits = PENetwork_15_io_to_pes_1_in_bits; // @[pe.scala 262:34]
  assign PE_45_io_data_0_in_valid = PENetwork_1_io_to_pes_4_in_valid; // @[pe.scala 262:34]
  assign PE_45_io_data_0_in_bits = PENetwork_1_io_to_pes_4_in_bits; // @[pe.scala 262:34]
  assign PE_46_clock = clock;
  assign PE_46_reset = reset;
  assign PE_46_io_data_2_in_valid = PENetwork_30_io_to_pes_2_in_valid; // @[pe.scala 262:34]
  assign PE_46_io_data_2_in_bits = PENetwork_30_io_to_pes_2_in_bits; // @[pe.scala 262:34]
  assign PE_46_io_data_2_sig_stat2trans = PENetwork_30_io_to_pes_2_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_46_io_data_2_out_ready = PENetwork_30_io_to_pes_2_out_ready; // @[pe.scala 268:49]
  assign PE_46_io_data_1_in_valid = PENetwork_15_io_to_pes_2_in_valid; // @[pe.scala 262:34]
  assign PE_46_io_data_1_in_bits = PENetwork_15_io_to_pes_2_in_bits; // @[pe.scala 262:34]
  assign PE_46_io_data_0_in_valid = PENetwork_2_io_to_pes_4_in_valid; // @[pe.scala 262:34]
  assign PE_46_io_data_0_in_bits = PENetwork_2_io_to_pes_4_in_bits; // @[pe.scala 262:34]
  assign PE_47_clock = clock;
  assign PE_47_reset = reset;
  assign PE_47_io_data_2_in_valid = PENetwork_30_io_to_pes_3_in_valid; // @[pe.scala 262:34]
  assign PE_47_io_data_2_in_bits = PENetwork_30_io_to_pes_3_in_bits; // @[pe.scala 262:34]
  assign PE_47_io_data_2_sig_stat2trans = PENetwork_30_io_to_pes_3_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_47_io_data_2_out_ready = PENetwork_30_io_to_pes_3_out_ready; // @[pe.scala 268:49]
  assign PE_47_io_data_1_in_valid = PENetwork_15_io_to_pes_3_in_valid; // @[pe.scala 262:34]
  assign PE_47_io_data_1_in_bits = PENetwork_15_io_to_pes_3_in_bits; // @[pe.scala 262:34]
  assign PE_47_io_data_0_in_valid = PENetwork_3_io_to_pes_4_in_valid; // @[pe.scala 262:34]
  assign PE_47_io_data_0_in_bits = PENetwork_3_io_to_pes_4_in_bits; // @[pe.scala 262:34]
  assign PE_48_clock = clock;
  assign PE_48_reset = reset;
  assign PE_48_io_data_2_in_valid = PENetwork_30_io_to_pes_4_in_valid; // @[pe.scala 262:34]
  assign PE_48_io_data_2_in_bits = PENetwork_30_io_to_pes_4_in_bits; // @[pe.scala 262:34]
  assign PE_48_io_data_2_sig_stat2trans = PENetwork_30_io_to_pes_4_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_48_io_data_2_out_ready = PENetwork_30_io_to_pes_4_out_ready; // @[pe.scala 268:49]
  assign PE_48_io_data_1_in_valid = PENetwork_15_io_to_pes_4_in_valid; // @[pe.scala 262:34]
  assign PE_48_io_data_1_in_bits = PENetwork_15_io_to_pes_4_in_bits; // @[pe.scala 262:34]
  assign PE_48_io_data_0_in_valid = PENetwork_4_io_to_pes_4_in_valid; // @[pe.scala 262:34]
  assign PE_48_io_data_0_in_bits = PENetwork_4_io_to_pes_4_in_bits; // @[pe.scala 262:34]
  assign PE_49_clock = clock;
  assign PE_49_reset = reset;
  assign PE_49_io_data_2_in_valid = PENetwork_30_io_to_pes_5_in_valid; // @[pe.scala 262:34]
  assign PE_49_io_data_2_in_bits = PENetwork_30_io_to_pes_5_in_bits; // @[pe.scala 262:34]
  assign PE_49_io_data_2_sig_stat2trans = PENetwork_30_io_to_pes_5_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_49_io_data_2_out_ready = PENetwork_30_io_to_pes_5_out_ready; // @[pe.scala 268:49]
  assign PE_49_io_data_1_in_valid = PENetwork_15_io_to_pes_5_in_valid; // @[pe.scala 262:34]
  assign PE_49_io_data_1_in_bits = PENetwork_15_io_to_pes_5_in_bits; // @[pe.scala 262:34]
  assign PE_49_io_data_0_in_valid = PENetwork_5_io_to_pes_4_in_valid; // @[pe.scala 262:34]
  assign PE_49_io_data_0_in_bits = PENetwork_5_io_to_pes_4_in_bits; // @[pe.scala 262:34]
  assign PE_50_clock = clock;
  assign PE_50_reset = reset;
  assign PE_50_io_data_2_in_valid = PENetwork_30_io_to_pes_6_in_valid; // @[pe.scala 262:34]
  assign PE_50_io_data_2_in_bits = PENetwork_30_io_to_pes_6_in_bits; // @[pe.scala 262:34]
  assign PE_50_io_data_2_sig_stat2trans = PENetwork_30_io_to_pes_6_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_50_io_data_2_out_ready = PENetwork_30_io_to_pes_6_out_ready; // @[pe.scala 268:49]
  assign PE_50_io_data_1_in_valid = PENetwork_15_io_to_pes_6_in_valid; // @[pe.scala 262:34]
  assign PE_50_io_data_1_in_bits = PENetwork_15_io_to_pes_6_in_bits; // @[pe.scala 262:34]
  assign PE_50_io_data_0_in_valid = PENetwork_6_io_to_pes_4_in_valid; // @[pe.scala 262:34]
  assign PE_50_io_data_0_in_bits = PENetwork_6_io_to_pes_4_in_bits; // @[pe.scala 262:34]
  assign PE_51_clock = clock;
  assign PE_51_reset = reset;
  assign PE_51_io_data_2_in_valid = PENetwork_30_io_to_pes_7_in_valid; // @[pe.scala 262:34]
  assign PE_51_io_data_2_in_bits = PENetwork_30_io_to_pes_7_in_bits; // @[pe.scala 262:34]
  assign PE_51_io_data_2_sig_stat2trans = PENetwork_30_io_to_pes_7_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_51_io_data_2_out_ready = PENetwork_30_io_to_pes_7_out_ready; // @[pe.scala 268:49]
  assign PE_51_io_data_1_in_valid = PENetwork_15_io_to_pes_7_in_valid; // @[pe.scala 262:34]
  assign PE_51_io_data_1_in_bits = PENetwork_15_io_to_pes_7_in_bits; // @[pe.scala 262:34]
  assign PE_51_io_data_0_in_valid = PENetwork_7_io_to_pes_4_in_valid; // @[pe.scala 262:34]
  assign PE_51_io_data_0_in_bits = PENetwork_7_io_to_pes_4_in_bits; // @[pe.scala 262:34]
  assign PE_52_clock = clock;
  assign PE_52_reset = reset;
  assign PE_52_io_data_2_in_valid = PENetwork_30_io_to_pes_8_in_valid; // @[pe.scala 262:34]
  assign PE_52_io_data_2_in_bits = PENetwork_30_io_to_pes_8_in_bits; // @[pe.scala 262:34]
  assign PE_52_io_data_2_sig_stat2trans = PENetwork_30_io_to_pes_8_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_52_io_data_2_out_ready = PENetwork_30_io_to_pes_8_out_ready; // @[pe.scala 268:49]
  assign PE_52_io_data_1_in_valid = PENetwork_15_io_to_pes_8_in_valid; // @[pe.scala 262:34]
  assign PE_52_io_data_1_in_bits = PENetwork_15_io_to_pes_8_in_bits; // @[pe.scala 262:34]
  assign PE_52_io_data_0_in_valid = PENetwork_8_io_to_pes_4_in_valid; // @[pe.scala 262:34]
  assign PE_52_io_data_0_in_bits = PENetwork_8_io_to_pes_4_in_bits; // @[pe.scala 262:34]
  assign PE_53_clock = clock;
  assign PE_53_reset = reset;
  assign PE_53_io_data_2_in_valid = PENetwork_30_io_to_pes_9_in_valid; // @[pe.scala 262:34]
  assign PE_53_io_data_2_in_bits = PENetwork_30_io_to_pes_9_in_bits; // @[pe.scala 262:34]
  assign PE_53_io_data_2_sig_stat2trans = PENetwork_30_io_to_pes_9_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_53_io_data_2_out_ready = PENetwork_30_io_to_pes_9_out_ready; // @[pe.scala 268:49]
  assign PE_53_io_data_1_in_valid = PENetwork_15_io_to_pes_9_in_valid; // @[pe.scala 262:34]
  assign PE_53_io_data_1_in_bits = PENetwork_15_io_to_pes_9_in_bits; // @[pe.scala 262:34]
  assign PE_53_io_data_0_in_valid = PENetwork_9_io_to_pes_4_in_valid; // @[pe.scala 262:34]
  assign PE_53_io_data_0_in_bits = PENetwork_9_io_to_pes_4_in_bits; // @[pe.scala 262:34]
  assign PE_54_clock = clock;
  assign PE_54_reset = reset;
  assign PE_54_io_data_2_in_valid = PENetwork_30_io_to_pes_10_in_valid; // @[pe.scala 262:34]
  assign PE_54_io_data_2_in_bits = PENetwork_30_io_to_pes_10_in_bits; // @[pe.scala 262:34]
  assign PE_54_io_data_2_sig_stat2trans = PENetwork_30_io_to_pes_10_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_54_io_data_2_out_ready = 1'h1; // @[pe.scala 268:49]
  assign PE_54_io_data_1_in_valid = PENetwork_15_io_to_pes_10_in_valid; // @[pe.scala 262:34]
  assign PE_54_io_data_1_in_bits = PENetwork_15_io_to_pes_10_in_bits; // @[pe.scala 262:34]
  assign PE_54_io_data_0_in_valid = PENetwork_10_io_to_pes_4_in_valid; // @[pe.scala 262:34]
  assign PE_54_io_data_0_in_bits = PENetwork_10_io_to_pes_4_in_bits; // @[pe.scala 262:34]
  assign PE_55_clock = clock;
  assign PE_55_reset = reset;
  assign PE_55_io_data_2_in_valid = 1'h0; // @[pe.scala 262:34]
  assign PE_55_io_data_2_in_bits = 256'h0; // @[pe.scala 262:34]
  assign PE_55_io_data_2_sig_stat2trans = PENetwork_31_io_to_pes_0_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_55_io_data_2_out_ready = PENetwork_31_io_to_pes_0_out_ready; // @[pe.scala 268:49]
  assign PE_55_io_data_1_in_valid = PENetwork_16_io_to_pes_0_in_valid; // @[pe.scala 262:34]
  assign PE_55_io_data_1_in_bits = PENetwork_16_io_to_pes_0_in_bits; // @[pe.scala 262:34]
  assign PE_55_io_data_0_in_valid = PENetwork_io_to_pes_5_in_valid; // @[pe.scala 262:34]
  assign PE_55_io_data_0_in_bits = PENetwork_io_to_pes_5_in_bits; // @[pe.scala 262:34]
  assign PE_56_clock = clock;
  assign PE_56_reset = reset;
  assign PE_56_io_data_2_in_valid = PENetwork_31_io_to_pes_1_in_valid; // @[pe.scala 262:34]
  assign PE_56_io_data_2_in_bits = PENetwork_31_io_to_pes_1_in_bits; // @[pe.scala 262:34]
  assign PE_56_io_data_2_sig_stat2trans = PENetwork_31_io_to_pes_1_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_56_io_data_2_out_ready = PENetwork_31_io_to_pes_1_out_ready; // @[pe.scala 268:49]
  assign PE_56_io_data_1_in_valid = PENetwork_16_io_to_pes_1_in_valid; // @[pe.scala 262:34]
  assign PE_56_io_data_1_in_bits = PENetwork_16_io_to_pes_1_in_bits; // @[pe.scala 262:34]
  assign PE_56_io_data_0_in_valid = PENetwork_1_io_to_pes_5_in_valid; // @[pe.scala 262:34]
  assign PE_56_io_data_0_in_bits = PENetwork_1_io_to_pes_5_in_bits; // @[pe.scala 262:34]
  assign PE_57_clock = clock;
  assign PE_57_reset = reset;
  assign PE_57_io_data_2_in_valid = PENetwork_31_io_to_pes_2_in_valid; // @[pe.scala 262:34]
  assign PE_57_io_data_2_in_bits = PENetwork_31_io_to_pes_2_in_bits; // @[pe.scala 262:34]
  assign PE_57_io_data_2_sig_stat2trans = PENetwork_31_io_to_pes_2_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_57_io_data_2_out_ready = PENetwork_31_io_to_pes_2_out_ready; // @[pe.scala 268:49]
  assign PE_57_io_data_1_in_valid = PENetwork_16_io_to_pes_2_in_valid; // @[pe.scala 262:34]
  assign PE_57_io_data_1_in_bits = PENetwork_16_io_to_pes_2_in_bits; // @[pe.scala 262:34]
  assign PE_57_io_data_0_in_valid = PENetwork_2_io_to_pes_5_in_valid; // @[pe.scala 262:34]
  assign PE_57_io_data_0_in_bits = PENetwork_2_io_to_pes_5_in_bits; // @[pe.scala 262:34]
  assign PE_58_clock = clock;
  assign PE_58_reset = reset;
  assign PE_58_io_data_2_in_valid = PENetwork_31_io_to_pes_3_in_valid; // @[pe.scala 262:34]
  assign PE_58_io_data_2_in_bits = PENetwork_31_io_to_pes_3_in_bits; // @[pe.scala 262:34]
  assign PE_58_io_data_2_sig_stat2trans = PENetwork_31_io_to_pes_3_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_58_io_data_2_out_ready = PENetwork_31_io_to_pes_3_out_ready; // @[pe.scala 268:49]
  assign PE_58_io_data_1_in_valid = PENetwork_16_io_to_pes_3_in_valid; // @[pe.scala 262:34]
  assign PE_58_io_data_1_in_bits = PENetwork_16_io_to_pes_3_in_bits; // @[pe.scala 262:34]
  assign PE_58_io_data_0_in_valid = PENetwork_3_io_to_pes_5_in_valid; // @[pe.scala 262:34]
  assign PE_58_io_data_0_in_bits = PENetwork_3_io_to_pes_5_in_bits; // @[pe.scala 262:34]
  assign PE_59_clock = clock;
  assign PE_59_reset = reset;
  assign PE_59_io_data_2_in_valid = PENetwork_31_io_to_pes_4_in_valid; // @[pe.scala 262:34]
  assign PE_59_io_data_2_in_bits = PENetwork_31_io_to_pes_4_in_bits; // @[pe.scala 262:34]
  assign PE_59_io_data_2_sig_stat2trans = PENetwork_31_io_to_pes_4_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_59_io_data_2_out_ready = PENetwork_31_io_to_pes_4_out_ready; // @[pe.scala 268:49]
  assign PE_59_io_data_1_in_valid = PENetwork_16_io_to_pes_4_in_valid; // @[pe.scala 262:34]
  assign PE_59_io_data_1_in_bits = PENetwork_16_io_to_pes_4_in_bits; // @[pe.scala 262:34]
  assign PE_59_io_data_0_in_valid = PENetwork_4_io_to_pes_5_in_valid; // @[pe.scala 262:34]
  assign PE_59_io_data_0_in_bits = PENetwork_4_io_to_pes_5_in_bits; // @[pe.scala 262:34]
  assign PE_60_clock = clock;
  assign PE_60_reset = reset;
  assign PE_60_io_data_2_in_valid = PENetwork_31_io_to_pes_5_in_valid; // @[pe.scala 262:34]
  assign PE_60_io_data_2_in_bits = PENetwork_31_io_to_pes_5_in_bits; // @[pe.scala 262:34]
  assign PE_60_io_data_2_sig_stat2trans = PENetwork_31_io_to_pes_5_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_60_io_data_2_out_ready = PENetwork_31_io_to_pes_5_out_ready; // @[pe.scala 268:49]
  assign PE_60_io_data_1_in_valid = PENetwork_16_io_to_pes_5_in_valid; // @[pe.scala 262:34]
  assign PE_60_io_data_1_in_bits = PENetwork_16_io_to_pes_5_in_bits; // @[pe.scala 262:34]
  assign PE_60_io_data_0_in_valid = PENetwork_5_io_to_pes_5_in_valid; // @[pe.scala 262:34]
  assign PE_60_io_data_0_in_bits = PENetwork_5_io_to_pes_5_in_bits; // @[pe.scala 262:34]
  assign PE_61_clock = clock;
  assign PE_61_reset = reset;
  assign PE_61_io_data_2_in_valid = PENetwork_31_io_to_pes_6_in_valid; // @[pe.scala 262:34]
  assign PE_61_io_data_2_in_bits = PENetwork_31_io_to_pes_6_in_bits; // @[pe.scala 262:34]
  assign PE_61_io_data_2_sig_stat2trans = PENetwork_31_io_to_pes_6_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_61_io_data_2_out_ready = PENetwork_31_io_to_pes_6_out_ready; // @[pe.scala 268:49]
  assign PE_61_io_data_1_in_valid = PENetwork_16_io_to_pes_6_in_valid; // @[pe.scala 262:34]
  assign PE_61_io_data_1_in_bits = PENetwork_16_io_to_pes_6_in_bits; // @[pe.scala 262:34]
  assign PE_61_io_data_0_in_valid = PENetwork_6_io_to_pes_5_in_valid; // @[pe.scala 262:34]
  assign PE_61_io_data_0_in_bits = PENetwork_6_io_to_pes_5_in_bits; // @[pe.scala 262:34]
  assign PE_62_clock = clock;
  assign PE_62_reset = reset;
  assign PE_62_io_data_2_in_valid = PENetwork_31_io_to_pes_7_in_valid; // @[pe.scala 262:34]
  assign PE_62_io_data_2_in_bits = PENetwork_31_io_to_pes_7_in_bits; // @[pe.scala 262:34]
  assign PE_62_io_data_2_sig_stat2trans = PENetwork_31_io_to_pes_7_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_62_io_data_2_out_ready = PENetwork_31_io_to_pes_7_out_ready; // @[pe.scala 268:49]
  assign PE_62_io_data_1_in_valid = PENetwork_16_io_to_pes_7_in_valid; // @[pe.scala 262:34]
  assign PE_62_io_data_1_in_bits = PENetwork_16_io_to_pes_7_in_bits; // @[pe.scala 262:34]
  assign PE_62_io_data_0_in_valid = PENetwork_7_io_to_pes_5_in_valid; // @[pe.scala 262:34]
  assign PE_62_io_data_0_in_bits = PENetwork_7_io_to_pes_5_in_bits; // @[pe.scala 262:34]
  assign PE_63_clock = clock;
  assign PE_63_reset = reset;
  assign PE_63_io_data_2_in_valid = PENetwork_31_io_to_pes_8_in_valid; // @[pe.scala 262:34]
  assign PE_63_io_data_2_in_bits = PENetwork_31_io_to_pes_8_in_bits; // @[pe.scala 262:34]
  assign PE_63_io_data_2_sig_stat2trans = PENetwork_31_io_to_pes_8_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_63_io_data_2_out_ready = PENetwork_31_io_to_pes_8_out_ready; // @[pe.scala 268:49]
  assign PE_63_io_data_1_in_valid = PENetwork_16_io_to_pes_8_in_valid; // @[pe.scala 262:34]
  assign PE_63_io_data_1_in_bits = PENetwork_16_io_to_pes_8_in_bits; // @[pe.scala 262:34]
  assign PE_63_io_data_0_in_valid = PENetwork_8_io_to_pes_5_in_valid; // @[pe.scala 262:34]
  assign PE_63_io_data_0_in_bits = PENetwork_8_io_to_pes_5_in_bits; // @[pe.scala 262:34]
  assign PE_64_clock = clock;
  assign PE_64_reset = reset;
  assign PE_64_io_data_2_in_valid = PENetwork_31_io_to_pes_9_in_valid; // @[pe.scala 262:34]
  assign PE_64_io_data_2_in_bits = PENetwork_31_io_to_pes_9_in_bits; // @[pe.scala 262:34]
  assign PE_64_io_data_2_sig_stat2trans = PENetwork_31_io_to_pes_9_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_64_io_data_2_out_ready = PENetwork_31_io_to_pes_9_out_ready; // @[pe.scala 268:49]
  assign PE_64_io_data_1_in_valid = PENetwork_16_io_to_pes_9_in_valid; // @[pe.scala 262:34]
  assign PE_64_io_data_1_in_bits = PENetwork_16_io_to_pes_9_in_bits; // @[pe.scala 262:34]
  assign PE_64_io_data_0_in_valid = PENetwork_9_io_to_pes_5_in_valid; // @[pe.scala 262:34]
  assign PE_64_io_data_0_in_bits = PENetwork_9_io_to_pes_5_in_bits; // @[pe.scala 262:34]
  assign PE_65_clock = clock;
  assign PE_65_reset = reset;
  assign PE_65_io_data_2_in_valid = PENetwork_31_io_to_pes_10_in_valid; // @[pe.scala 262:34]
  assign PE_65_io_data_2_in_bits = PENetwork_31_io_to_pes_10_in_bits; // @[pe.scala 262:34]
  assign PE_65_io_data_2_sig_stat2trans = PENetwork_31_io_to_pes_10_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_65_io_data_2_out_ready = 1'h1; // @[pe.scala 268:49]
  assign PE_65_io_data_1_in_valid = PENetwork_16_io_to_pes_10_in_valid; // @[pe.scala 262:34]
  assign PE_65_io_data_1_in_bits = PENetwork_16_io_to_pes_10_in_bits; // @[pe.scala 262:34]
  assign PE_65_io_data_0_in_valid = PENetwork_10_io_to_pes_5_in_valid; // @[pe.scala 262:34]
  assign PE_65_io_data_0_in_bits = PENetwork_10_io_to_pes_5_in_bits; // @[pe.scala 262:34]
  assign PE_66_clock = clock;
  assign PE_66_reset = reset;
  assign PE_66_io_data_2_in_valid = 1'h0; // @[pe.scala 262:34]
  assign PE_66_io_data_2_in_bits = 256'h0; // @[pe.scala 262:34]
  assign PE_66_io_data_2_sig_stat2trans = PENetwork_32_io_to_pes_0_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_66_io_data_2_out_ready = PENetwork_32_io_to_pes_0_out_ready; // @[pe.scala 268:49]
  assign PE_66_io_data_1_in_valid = PENetwork_17_io_to_pes_0_in_valid; // @[pe.scala 262:34]
  assign PE_66_io_data_1_in_bits = PENetwork_17_io_to_pes_0_in_bits; // @[pe.scala 262:34]
  assign PE_66_io_data_0_in_valid = PENetwork_io_to_pes_6_in_valid; // @[pe.scala 262:34]
  assign PE_66_io_data_0_in_bits = PENetwork_io_to_pes_6_in_bits; // @[pe.scala 262:34]
  assign PE_67_clock = clock;
  assign PE_67_reset = reset;
  assign PE_67_io_data_2_in_valid = PENetwork_32_io_to_pes_1_in_valid; // @[pe.scala 262:34]
  assign PE_67_io_data_2_in_bits = PENetwork_32_io_to_pes_1_in_bits; // @[pe.scala 262:34]
  assign PE_67_io_data_2_sig_stat2trans = PENetwork_32_io_to_pes_1_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_67_io_data_2_out_ready = PENetwork_32_io_to_pes_1_out_ready; // @[pe.scala 268:49]
  assign PE_67_io_data_1_in_valid = PENetwork_17_io_to_pes_1_in_valid; // @[pe.scala 262:34]
  assign PE_67_io_data_1_in_bits = PENetwork_17_io_to_pes_1_in_bits; // @[pe.scala 262:34]
  assign PE_67_io_data_0_in_valid = PENetwork_1_io_to_pes_6_in_valid; // @[pe.scala 262:34]
  assign PE_67_io_data_0_in_bits = PENetwork_1_io_to_pes_6_in_bits; // @[pe.scala 262:34]
  assign PE_68_clock = clock;
  assign PE_68_reset = reset;
  assign PE_68_io_data_2_in_valid = PENetwork_32_io_to_pes_2_in_valid; // @[pe.scala 262:34]
  assign PE_68_io_data_2_in_bits = PENetwork_32_io_to_pes_2_in_bits; // @[pe.scala 262:34]
  assign PE_68_io_data_2_sig_stat2trans = PENetwork_32_io_to_pes_2_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_68_io_data_2_out_ready = PENetwork_32_io_to_pes_2_out_ready; // @[pe.scala 268:49]
  assign PE_68_io_data_1_in_valid = PENetwork_17_io_to_pes_2_in_valid; // @[pe.scala 262:34]
  assign PE_68_io_data_1_in_bits = PENetwork_17_io_to_pes_2_in_bits; // @[pe.scala 262:34]
  assign PE_68_io_data_0_in_valid = PENetwork_2_io_to_pes_6_in_valid; // @[pe.scala 262:34]
  assign PE_68_io_data_0_in_bits = PENetwork_2_io_to_pes_6_in_bits; // @[pe.scala 262:34]
  assign PE_69_clock = clock;
  assign PE_69_reset = reset;
  assign PE_69_io_data_2_in_valid = PENetwork_32_io_to_pes_3_in_valid; // @[pe.scala 262:34]
  assign PE_69_io_data_2_in_bits = PENetwork_32_io_to_pes_3_in_bits; // @[pe.scala 262:34]
  assign PE_69_io_data_2_sig_stat2trans = PENetwork_32_io_to_pes_3_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_69_io_data_2_out_ready = PENetwork_32_io_to_pes_3_out_ready; // @[pe.scala 268:49]
  assign PE_69_io_data_1_in_valid = PENetwork_17_io_to_pes_3_in_valid; // @[pe.scala 262:34]
  assign PE_69_io_data_1_in_bits = PENetwork_17_io_to_pes_3_in_bits; // @[pe.scala 262:34]
  assign PE_69_io_data_0_in_valid = PENetwork_3_io_to_pes_6_in_valid; // @[pe.scala 262:34]
  assign PE_69_io_data_0_in_bits = PENetwork_3_io_to_pes_6_in_bits; // @[pe.scala 262:34]
  assign PE_70_clock = clock;
  assign PE_70_reset = reset;
  assign PE_70_io_data_2_in_valid = PENetwork_32_io_to_pes_4_in_valid; // @[pe.scala 262:34]
  assign PE_70_io_data_2_in_bits = PENetwork_32_io_to_pes_4_in_bits; // @[pe.scala 262:34]
  assign PE_70_io_data_2_sig_stat2trans = PENetwork_32_io_to_pes_4_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_70_io_data_2_out_ready = PENetwork_32_io_to_pes_4_out_ready; // @[pe.scala 268:49]
  assign PE_70_io_data_1_in_valid = PENetwork_17_io_to_pes_4_in_valid; // @[pe.scala 262:34]
  assign PE_70_io_data_1_in_bits = PENetwork_17_io_to_pes_4_in_bits; // @[pe.scala 262:34]
  assign PE_70_io_data_0_in_valid = PENetwork_4_io_to_pes_6_in_valid; // @[pe.scala 262:34]
  assign PE_70_io_data_0_in_bits = PENetwork_4_io_to_pes_6_in_bits; // @[pe.scala 262:34]
  assign PE_71_clock = clock;
  assign PE_71_reset = reset;
  assign PE_71_io_data_2_in_valid = PENetwork_32_io_to_pes_5_in_valid; // @[pe.scala 262:34]
  assign PE_71_io_data_2_in_bits = PENetwork_32_io_to_pes_5_in_bits; // @[pe.scala 262:34]
  assign PE_71_io_data_2_sig_stat2trans = PENetwork_32_io_to_pes_5_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_71_io_data_2_out_ready = PENetwork_32_io_to_pes_5_out_ready; // @[pe.scala 268:49]
  assign PE_71_io_data_1_in_valid = PENetwork_17_io_to_pes_5_in_valid; // @[pe.scala 262:34]
  assign PE_71_io_data_1_in_bits = PENetwork_17_io_to_pes_5_in_bits; // @[pe.scala 262:34]
  assign PE_71_io_data_0_in_valid = PENetwork_5_io_to_pes_6_in_valid; // @[pe.scala 262:34]
  assign PE_71_io_data_0_in_bits = PENetwork_5_io_to_pes_6_in_bits; // @[pe.scala 262:34]
  assign PE_72_clock = clock;
  assign PE_72_reset = reset;
  assign PE_72_io_data_2_in_valid = PENetwork_32_io_to_pes_6_in_valid; // @[pe.scala 262:34]
  assign PE_72_io_data_2_in_bits = PENetwork_32_io_to_pes_6_in_bits; // @[pe.scala 262:34]
  assign PE_72_io_data_2_sig_stat2trans = PENetwork_32_io_to_pes_6_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_72_io_data_2_out_ready = PENetwork_32_io_to_pes_6_out_ready; // @[pe.scala 268:49]
  assign PE_72_io_data_1_in_valid = PENetwork_17_io_to_pes_6_in_valid; // @[pe.scala 262:34]
  assign PE_72_io_data_1_in_bits = PENetwork_17_io_to_pes_6_in_bits; // @[pe.scala 262:34]
  assign PE_72_io_data_0_in_valid = PENetwork_6_io_to_pes_6_in_valid; // @[pe.scala 262:34]
  assign PE_72_io_data_0_in_bits = PENetwork_6_io_to_pes_6_in_bits; // @[pe.scala 262:34]
  assign PE_73_clock = clock;
  assign PE_73_reset = reset;
  assign PE_73_io_data_2_in_valid = PENetwork_32_io_to_pes_7_in_valid; // @[pe.scala 262:34]
  assign PE_73_io_data_2_in_bits = PENetwork_32_io_to_pes_7_in_bits; // @[pe.scala 262:34]
  assign PE_73_io_data_2_sig_stat2trans = PENetwork_32_io_to_pes_7_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_73_io_data_2_out_ready = PENetwork_32_io_to_pes_7_out_ready; // @[pe.scala 268:49]
  assign PE_73_io_data_1_in_valid = PENetwork_17_io_to_pes_7_in_valid; // @[pe.scala 262:34]
  assign PE_73_io_data_1_in_bits = PENetwork_17_io_to_pes_7_in_bits; // @[pe.scala 262:34]
  assign PE_73_io_data_0_in_valid = PENetwork_7_io_to_pes_6_in_valid; // @[pe.scala 262:34]
  assign PE_73_io_data_0_in_bits = PENetwork_7_io_to_pes_6_in_bits; // @[pe.scala 262:34]
  assign PE_74_clock = clock;
  assign PE_74_reset = reset;
  assign PE_74_io_data_2_in_valid = PENetwork_32_io_to_pes_8_in_valid; // @[pe.scala 262:34]
  assign PE_74_io_data_2_in_bits = PENetwork_32_io_to_pes_8_in_bits; // @[pe.scala 262:34]
  assign PE_74_io_data_2_sig_stat2trans = PENetwork_32_io_to_pes_8_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_74_io_data_2_out_ready = PENetwork_32_io_to_pes_8_out_ready; // @[pe.scala 268:49]
  assign PE_74_io_data_1_in_valid = PENetwork_17_io_to_pes_8_in_valid; // @[pe.scala 262:34]
  assign PE_74_io_data_1_in_bits = PENetwork_17_io_to_pes_8_in_bits; // @[pe.scala 262:34]
  assign PE_74_io_data_0_in_valid = PENetwork_8_io_to_pes_6_in_valid; // @[pe.scala 262:34]
  assign PE_74_io_data_0_in_bits = PENetwork_8_io_to_pes_6_in_bits; // @[pe.scala 262:34]
  assign PE_75_clock = clock;
  assign PE_75_reset = reset;
  assign PE_75_io_data_2_in_valid = PENetwork_32_io_to_pes_9_in_valid; // @[pe.scala 262:34]
  assign PE_75_io_data_2_in_bits = PENetwork_32_io_to_pes_9_in_bits; // @[pe.scala 262:34]
  assign PE_75_io_data_2_sig_stat2trans = PENetwork_32_io_to_pes_9_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_75_io_data_2_out_ready = PENetwork_32_io_to_pes_9_out_ready; // @[pe.scala 268:49]
  assign PE_75_io_data_1_in_valid = PENetwork_17_io_to_pes_9_in_valid; // @[pe.scala 262:34]
  assign PE_75_io_data_1_in_bits = PENetwork_17_io_to_pes_9_in_bits; // @[pe.scala 262:34]
  assign PE_75_io_data_0_in_valid = PENetwork_9_io_to_pes_6_in_valid; // @[pe.scala 262:34]
  assign PE_75_io_data_0_in_bits = PENetwork_9_io_to_pes_6_in_bits; // @[pe.scala 262:34]
  assign PE_76_clock = clock;
  assign PE_76_reset = reset;
  assign PE_76_io_data_2_in_valid = PENetwork_32_io_to_pes_10_in_valid; // @[pe.scala 262:34]
  assign PE_76_io_data_2_in_bits = PENetwork_32_io_to_pes_10_in_bits; // @[pe.scala 262:34]
  assign PE_76_io_data_2_sig_stat2trans = PENetwork_32_io_to_pes_10_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_76_io_data_2_out_ready = 1'h1; // @[pe.scala 268:49]
  assign PE_76_io_data_1_in_valid = PENetwork_17_io_to_pes_10_in_valid; // @[pe.scala 262:34]
  assign PE_76_io_data_1_in_bits = PENetwork_17_io_to_pes_10_in_bits; // @[pe.scala 262:34]
  assign PE_76_io_data_0_in_valid = PENetwork_10_io_to_pes_6_in_valid; // @[pe.scala 262:34]
  assign PE_76_io_data_0_in_bits = PENetwork_10_io_to_pes_6_in_bits; // @[pe.scala 262:34]
  assign PE_77_clock = clock;
  assign PE_77_reset = reset;
  assign PE_77_io_data_2_in_valid = 1'h0; // @[pe.scala 262:34]
  assign PE_77_io_data_2_in_bits = 256'h0; // @[pe.scala 262:34]
  assign PE_77_io_data_2_sig_stat2trans = PENetwork_33_io_to_pes_0_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_77_io_data_2_out_ready = PENetwork_33_io_to_pes_0_out_ready; // @[pe.scala 268:49]
  assign PE_77_io_data_1_in_valid = PENetwork_18_io_to_pes_0_in_valid; // @[pe.scala 262:34]
  assign PE_77_io_data_1_in_bits = PENetwork_18_io_to_pes_0_in_bits; // @[pe.scala 262:34]
  assign PE_77_io_data_0_in_valid = PENetwork_io_to_pes_7_in_valid; // @[pe.scala 262:34]
  assign PE_77_io_data_0_in_bits = PENetwork_io_to_pes_7_in_bits; // @[pe.scala 262:34]
  assign PE_78_clock = clock;
  assign PE_78_reset = reset;
  assign PE_78_io_data_2_in_valid = PENetwork_33_io_to_pes_1_in_valid; // @[pe.scala 262:34]
  assign PE_78_io_data_2_in_bits = PENetwork_33_io_to_pes_1_in_bits; // @[pe.scala 262:34]
  assign PE_78_io_data_2_sig_stat2trans = PENetwork_33_io_to_pes_1_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_78_io_data_2_out_ready = PENetwork_33_io_to_pes_1_out_ready; // @[pe.scala 268:49]
  assign PE_78_io_data_1_in_valid = PENetwork_18_io_to_pes_1_in_valid; // @[pe.scala 262:34]
  assign PE_78_io_data_1_in_bits = PENetwork_18_io_to_pes_1_in_bits; // @[pe.scala 262:34]
  assign PE_78_io_data_0_in_valid = PENetwork_1_io_to_pes_7_in_valid; // @[pe.scala 262:34]
  assign PE_78_io_data_0_in_bits = PENetwork_1_io_to_pes_7_in_bits; // @[pe.scala 262:34]
  assign PE_79_clock = clock;
  assign PE_79_reset = reset;
  assign PE_79_io_data_2_in_valid = PENetwork_33_io_to_pes_2_in_valid; // @[pe.scala 262:34]
  assign PE_79_io_data_2_in_bits = PENetwork_33_io_to_pes_2_in_bits; // @[pe.scala 262:34]
  assign PE_79_io_data_2_sig_stat2trans = PENetwork_33_io_to_pes_2_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_79_io_data_2_out_ready = PENetwork_33_io_to_pes_2_out_ready; // @[pe.scala 268:49]
  assign PE_79_io_data_1_in_valid = PENetwork_18_io_to_pes_2_in_valid; // @[pe.scala 262:34]
  assign PE_79_io_data_1_in_bits = PENetwork_18_io_to_pes_2_in_bits; // @[pe.scala 262:34]
  assign PE_79_io_data_0_in_valid = PENetwork_2_io_to_pes_7_in_valid; // @[pe.scala 262:34]
  assign PE_79_io_data_0_in_bits = PENetwork_2_io_to_pes_7_in_bits; // @[pe.scala 262:34]
  assign PE_80_clock = clock;
  assign PE_80_reset = reset;
  assign PE_80_io_data_2_in_valid = PENetwork_33_io_to_pes_3_in_valid; // @[pe.scala 262:34]
  assign PE_80_io_data_2_in_bits = PENetwork_33_io_to_pes_3_in_bits; // @[pe.scala 262:34]
  assign PE_80_io_data_2_sig_stat2trans = PENetwork_33_io_to_pes_3_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_80_io_data_2_out_ready = PENetwork_33_io_to_pes_3_out_ready; // @[pe.scala 268:49]
  assign PE_80_io_data_1_in_valid = PENetwork_18_io_to_pes_3_in_valid; // @[pe.scala 262:34]
  assign PE_80_io_data_1_in_bits = PENetwork_18_io_to_pes_3_in_bits; // @[pe.scala 262:34]
  assign PE_80_io_data_0_in_valid = PENetwork_3_io_to_pes_7_in_valid; // @[pe.scala 262:34]
  assign PE_80_io_data_0_in_bits = PENetwork_3_io_to_pes_7_in_bits; // @[pe.scala 262:34]
  assign PE_81_clock = clock;
  assign PE_81_reset = reset;
  assign PE_81_io_data_2_in_valid = PENetwork_33_io_to_pes_4_in_valid; // @[pe.scala 262:34]
  assign PE_81_io_data_2_in_bits = PENetwork_33_io_to_pes_4_in_bits; // @[pe.scala 262:34]
  assign PE_81_io_data_2_sig_stat2trans = PENetwork_33_io_to_pes_4_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_81_io_data_2_out_ready = PENetwork_33_io_to_pes_4_out_ready; // @[pe.scala 268:49]
  assign PE_81_io_data_1_in_valid = PENetwork_18_io_to_pes_4_in_valid; // @[pe.scala 262:34]
  assign PE_81_io_data_1_in_bits = PENetwork_18_io_to_pes_4_in_bits; // @[pe.scala 262:34]
  assign PE_81_io_data_0_in_valid = PENetwork_4_io_to_pes_7_in_valid; // @[pe.scala 262:34]
  assign PE_81_io_data_0_in_bits = PENetwork_4_io_to_pes_7_in_bits; // @[pe.scala 262:34]
  assign PE_82_clock = clock;
  assign PE_82_reset = reset;
  assign PE_82_io_data_2_in_valid = PENetwork_33_io_to_pes_5_in_valid; // @[pe.scala 262:34]
  assign PE_82_io_data_2_in_bits = PENetwork_33_io_to_pes_5_in_bits; // @[pe.scala 262:34]
  assign PE_82_io_data_2_sig_stat2trans = PENetwork_33_io_to_pes_5_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_82_io_data_2_out_ready = PENetwork_33_io_to_pes_5_out_ready; // @[pe.scala 268:49]
  assign PE_82_io_data_1_in_valid = PENetwork_18_io_to_pes_5_in_valid; // @[pe.scala 262:34]
  assign PE_82_io_data_1_in_bits = PENetwork_18_io_to_pes_5_in_bits; // @[pe.scala 262:34]
  assign PE_82_io_data_0_in_valid = PENetwork_5_io_to_pes_7_in_valid; // @[pe.scala 262:34]
  assign PE_82_io_data_0_in_bits = PENetwork_5_io_to_pes_7_in_bits; // @[pe.scala 262:34]
  assign PE_83_clock = clock;
  assign PE_83_reset = reset;
  assign PE_83_io_data_2_in_valid = PENetwork_33_io_to_pes_6_in_valid; // @[pe.scala 262:34]
  assign PE_83_io_data_2_in_bits = PENetwork_33_io_to_pes_6_in_bits; // @[pe.scala 262:34]
  assign PE_83_io_data_2_sig_stat2trans = PENetwork_33_io_to_pes_6_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_83_io_data_2_out_ready = PENetwork_33_io_to_pes_6_out_ready; // @[pe.scala 268:49]
  assign PE_83_io_data_1_in_valid = PENetwork_18_io_to_pes_6_in_valid; // @[pe.scala 262:34]
  assign PE_83_io_data_1_in_bits = PENetwork_18_io_to_pes_6_in_bits; // @[pe.scala 262:34]
  assign PE_83_io_data_0_in_valid = PENetwork_6_io_to_pes_7_in_valid; // @[pe.scala 262:34]
  assign PE_83_io_data_0_in_bits = PENetwork_6_io_to_pes_7_in_bits; // @[pe.scala 262:34]
  assign PE_84_clock = clock;
  assign PE_84_reset = reset;
  assign PE_84_io_data_2_in_valid = PENetwork_33_io_to_pes_7_in_valid; // @[pe.scala 262:34]
  assign PE_84_io_data_2_in_bits = PENetwork_33_io_to_pes_7_in_bits; // @[pe.scala 262:34]
  assign PE_84_io_data_2_sig_stat2trans = PENetwork_33_io_to_pes_7_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_84_io_data_2_out_ready = PENetwork_33_io_to_pes_7_out_ready; // @[pe.scala 268:49]
  assign PE_84_io_data_1_in_valid = PENetwork_18_io_to_pes_7_in_valid; // @[pe.scala 262:34]
  assign PE_84_io_data_1_in_bits = PENetwork_18_io_to_pes_7_in_bits; // @[pe.scala 262:34]
  assign PE_84_io_data_0_in_valid = PENetwork_7_io_to_pes_7_in_valid; // @[pe.scala 262:34]
  assign PE_84_io_data_0_in_bits = PENetwork_7_io_to_pes_7_in_bits; // @[pe.scala 262:34]
  assign PE_85_clock = clock;
  assign PE_85_reset = reset;
  assign PE_85_io_data_2_in_valid = PENetwork_33_io_to_pes_8_in_valid; // @[pe.scala 262:34]
  assign PE_85_io_data_2_in_bits = PENetwork_33_io_to_pes_8_in_bits; // @[pe.scala 262:34]
  assign PE_85_io_data_2_sig_stat2trans = PENetwork_33_io_to_pes_8_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_85_io_data_2_out_ready = PENetwork_33_io_to_pes_8_out_ready; // @[pe.scala 268:49]
  assign PE_85_io_data_1_in_valid = PENetwork_18_io_to_pes_8_in_valid; // @[pe.scala 262:34]
  assign PE_85_io_data_1_in_bits = PENetwork_18_io_to_pes_8_in_bits; // @[pe.scala 262:34]
  assign PE_85_io_data_0_in_valid = PENetwork_8_io_to_pes_7_in_valid; // @[pe.scala 262:34]
  assign PE_85_io_data_0_in_bits = PENetwork_8_io_to_pes_7_in_bits; // @[pe.scala 262:34]
  assign PE_86_clock = clock;
  assign PE_86_reset = reset;
  assign PE_86_io_data_2_in_valid = PENetwork_33_io_to_pes_9_in_valid; // @[pe.scala 262:34]
  assign PE_86_io_data_2_in_bits = PENetwork_33_io_to_pes_9_in_bits; // @[pe.scala 262:34]
  assign PE_86_io_data_2_sig_stat2trans = PENetwork_33_io_to_pes_9_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_86_io_data_2_out_ready = PENetwork_33_io_to_pes_9_out_ready; // @[pe.scala 268:49]
  assign PE_86_io_data_1_in_valid = PENetwork_18_io_to_pes_9_in_valid; // @[pe.scala 262:34]
  assign PE_86_io_data_1_in_bits = PENetwork_18_io_to_pes_9_in_bits; // @[pe.scala 262:34]
  assign PE_86_io_data_0_in_valid = PENetwork_9_io_to_pes_7_in_valid; // @[pe.scala 262:34]
  assign PE_86_io_data_0_in_bits = PENetwork_9_io_to_pes_7_in_bits; // @[pe.scala 262:34]
  assign PE_87_clock = clock;
  assign PE_87_reset = reset;
  assign PE_87_io_data_2_in_valid = PENetwork_33_io_to_pes_10_in_valid; // @[pe.scala 262:34]
  assign PE_87_io_data_2_in_bits = PENetwork_33_io_to_pes_10_in_bits; // @[pe.scala 262:34]
  assign PE_87_io_data_2_sig_stat2trans = PENetwork_33_io_to_pes_10_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_87_io_data_2_out_ready = 1'h1; // @[pe.scala 268:49]
  assign PE_87_io_data_1_in_valid = PENetwork_18_io_to_pes_10_in_valid; // @[pe.scala 262:34]
  assign PE_87_io_data_1_in_bits = PENetwork_18_io_to_pes_10_in_bits; // @[pe.scala 262:34]
  assign PE_87_io_data_0_in_valid = PENetwork_10_io_to_pes_7_in_valid; // @[pe.scala 262:34]
  assign PE_87_io_data_0_in_bits = PENetwork_10_io_to_pes_7_in_bits; // @[pe.scala 262:34]
  assign PE_88_clock = clock;
  assign PE_88_reset = reset;
  assign PE_88_io_data_2_in_valid = 1'h0; // @[pe.scala 262:34]
  assign PE_88_io_data_2_in_bits = 256'h0; // @[pe.scala 262:34]
  assign PE_88_io_data_2_sig_stat2trans = PENetwork_34_io_to_pes_0_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_88_io_data_2_out_ready = PENetwork_34_io_to_pes_0_out_ready; // @[pe.scala 268:49]
  assign PE_88_io_data_1_in_valid = PENetwork_19_io_to_pes_0_in_valid; // @[pe.scala 262:34]
  assign PE_88_io_data_1_in_bits = PENetwork_19_io_to_pes_0_in_bits; // @[pe.scala 262:34]
  assign PE_88_io_data_0_in_valid = PENetwork_io_to_pes_8_in_valid; // @[pe.scala 262:34]
  assign PE_88_io_data_0_in_bits = PENetwork_io_to_pes_8_in_bits; // @[pe.scala 262:34]
  assign PE_89_clock = clock;
  assign PE_89_reset = reset;
  assign PE_89_io_data_2_in_valid = PENetwork_34_io_to_pes_1_in_valid; // @[pe.scala 262:34]
  assign PE_89_io_data_2_in_bits = PENetwork_34_io_to_pes_1_in_bits; // @[pe.scala 262:34]
  assign PE_89_io_data_2_sig_stat2trans = PENetwork_34_io_to_pes_1_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_89_io_data_2_out_ready = PENetwork_34_io_to_pes_1_out_ready; // @[pe.scala 268:49]
  assign PE_89_io_data_1_in_valid = PENetwork_19_io_to_pes_1_in_valid; // @[pe.scala 262:34]
  assign PE_89_io_data_1_in_bits = PENetwork_19_io_to_pes_1_in_bits; // @[pe.scala 262:34]
  assign PE_89_io_data_0_in_valid = PENetwork_1_io_to_pes_8_in_valid; // @[pe.scala 262:34]
  assign PE_89_io_data_0_in_bits = PENetwork_1_io_to_pes_8_in_bits; // @[pe.scala 262:34]
  assign PE_90_clock = clock;
  assign PE_90_reset = reset;
  assign PE_90_io_data_2_in_valid = PENetwork_34_io_to_pes_2_in_valid; // @[pe.scala 262:34]
  assign PE_90_io_data_2_in_bits = PENetwork_34_io_to_pes_2_in_bits; // @[pe.scala 262:34]
  assign PE_90_io_data_2_sig_stat2trans = PENetwork_34_io_to_pes_2_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_90_io_data_2_out_ready = PENetwork_34_io_to_pes_2_out_ready; // @[pe.scala 268:49]
  assign PE_90_io_data_1_in_valid = PENetwork_19_io_to_pes_2_in_valid; // @[pe.scala 262:34]
  assign PE_90_io_data_1_in_bits = PENetwork_19_io_to_pes_2_in_bits; // @[pe.scala 262:34]
  assign PE_90_io_data_0_in_valid = PENetwork_2_io_to_pes_8_in_valid; // @[pe.scala 262:34]
  assign PE_90_io_data_0_in_bits = PENetwork_2_io_to_pes_8_in_bits; // @[pe.scala 262:34]
  assign PE_91_clock = clock;
  assign PE_91_reset = reset;
  assign PE_91_io_data_2_in_valid = PENetwork_34_io_to_pes_3_in_valid; // @[pe.scala 262:34]
  assign PE_91_io_data_2_in_bits = PENetwork_34_io_to_pes_3_in_bits; // @[pe.scala 262:34]
  assign PE_91_io_data_2_sig_stat2trans = PENetwork_34_io_to_pes_3_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_91_io_data_2_out_ready = PENetwork_34_io_to_pes_3_out_ready; // @[pe.scala 268:49]
  assign PE_91_io_data_1_in_valid = PENetwork_19_io_to_pes_3_in_valid; // @[pe.scala 262:34]
  assign PE_91_io_data_1_in_bits = PENetwork_19_io_to_pes_3_in_bits; // @[pe.scala 262:34]
  assign PE_91_io_data_0_in_valid = PENetwork_3_io_to_pes_8_in_valid; // @[pe.scala 262:34]
  assign PE_91_io_data_0_in_bits = PENetwork_3_io_to_pes_8_in_bits; // @[pe.scala 262:34]
  assign PE_92_clock = clock;
  assign PE_92_reset = reset;
  assign PE_92_io_data_2_in_valid = PENetwork_34_io_to_pes_4_in_valid; // @[pe.scala 262:34]
  assign PE_92_io_data_2_in_bits = PENetwork_34_io_to_pes_4_in_bits; // @[pe.scala 262:34]
  assign PE_92_io_data_2_sig_stat2trans = PENetwork_34_io_to_pes_4_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_92_io_data_2_out_ready = PENetwork_34_io_to_pes_4_out_ready; // @[pe.scala 268:49]
  assign PE_92_io_data_1_in_valid = PENetwork_19_io_to_pes_4_in_valid; // @[pe.scala 262:34]
  assign PE_92_io_data_1_in_bits = PENetwork_19_io_to_pes_4_in_bits; // @[pe.scala 262:34]
  assign PE_92_io_data_0_in_valid = PENetwork_4_io_to_pes_8_in_valid; // @[pe.scala 262:34]
  assign PE_92_io_data_0_in_bits = PENetwork_4_io_to_pes_8_in_bits; // @[pe.scala 262:34]
  assign PE_93_clock = clock;
  assign PE_93_reset = reset;
  assign PE_93_io_data_2_in_valid = PENetwork_34_io_to_pes_5_in_valid; // @[pe.scala 262:34]
  assign PE_93_io_data_2_in_bits = PENetwork_34_io_to_pes_5_in_bits; // @[pe.scala 262:34]
  assign PE_93_io_data_2_sig_stat2trans = PENetwork_34_io_to_pes_5_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_93_io_data_2_out_ready = PENetwork_34_io_to_pes_5_out_ready; // @[pe.scala 268:49]
  assign PE_93_io_data_1_in_valid = PENetwork_19_io_to_pes_5_in_valid; // @[pe.scala 262:34]
  assign PE_93_io_data_1_in_bits = PENetwork_19_io_to_pes_5_in_bits; // @[pe.scala 262:34]
  assign PE_93_io_data_0_in_valid = PENetwork_5_io_to_pes_8_in_valid; // @[pe.scala 262:34]
  assign PE_93_io_data_0_in_bits = PENetwork_5_io_to_pes_8_in_bits; // @[pe.scala 262:34]
  assign PE_94_clock = clock;
  assign PE_94_reset = reset;
  assign PE_94_io_data_2_in_valid = PENetwork_34_io_to_pes_6_in_valid; // @[pe.scala 262:34]
  assign PE_94_io_data_2_in_bits = PENetwork_34_io_to_pes_6_in_bits; // @[pe.scala 262:34]
  assign PE_94_io_data_2_sig_stat2trans = PENetwork_34_io_to_pes_6_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_94_io_data_2_out_ready = PENetwork_34_io_to_pes_6_out_ready; // @[pe.scala 268:49]
  assign PE_94_io_data_1_in_valid = PENetwork_19_io_to_pes_6_in_valid; // @[pe.scala 262:34]
  assign PE_94_io_data_1_in_bits = PENetwork_19_io_to_pes_6_in_bits; // @[pe.scala 262:34]
  assign PE_94_io_data_0_in_valid = PENetwork_6_io_to_pes_8_in_valid; // @[pe.scala 262:34]
  assign PE_94_io_data_0_in_bits = PENetwork_6_io_to_pes_8_in_bits; // @[pe.scala 262:34]
  assign PE_95_clock = clock;
  assign PE_95_reset = reset;
  assign PE_95_io_data_2_in_valid = PENetwork_34_io_to_pes_7_in_valid; // @[pe.scala 262:34]
  assign PE_95_io_data_2_in_bits = PENetwork_34_io_to_pes_7_in_bits; // @[pe.scala 262:34]
  assign PE_95_io_data_2_sig_stat2trans = PENetwork_34_io_to_pes_7_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_95_io_data_2_out_ready = PENetwork_34_io_to_pes_7_out_ready; // @[pe.scala 268:49]
  assign PE_95_io_data_1_in_valid = PENetwork_19_io_to_pes_7_in_valid; // @[pe.scala 262:34]
  assign PE_95_io_data_1_in_bits = PENetwork_19_io_to_pes_7_in_bits; // @[pe.scala 262:34]
  assign PE_95_io_data_0_in_valid = PENetwork_7_io_to_pes_8_in_valid; // @[pe.scala 262:34]
  assign PE_95_io_data_0_in_bits = PENetwork_7_io_to_pes_8_in_bits; // @[pe.scala 262:34]
  assign PE_96_clock = clock;
  assign PE_96_reset = reset;
  assign PE_96_io_data_2_in_valid = PENetwork_34_io_to_pes_8_in_valid; // @[pe.scala 262:34]
  assign PE_96_io_data_2_in_bits = PENetwork_34_io_to_pes_8_in_bits; // @[pe.scala 262:34]
  assign PE_96_io_data_2_sig_stat2trans = PENetwork_34_io_to_pes_8_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_96_io_data_2_out_ready = PENetwork_34_io_to_pes_8_out_ready; // @[pe.scala 268:49]
  assign PE_96_io_data_1_in_valid = PENetwork_19_io_to_pes_8_in_valid; // @[pe.scala 262:34]
  assign PE_96_io_data_1_in_bits = PENetwork_19_io_to_pes_8_in_bits; // @[pe.scala 262:34]
  assign PE_96_io_data_0_in_valid = PENetwork_8_io_to_pes_8_in_valid; // @[pe.scala 262:34]
  assign PE_96_io_data_0_in_bits = PENetwork_8_io_to_pes_8_in_bits; // @[pe.scala 262:34]
  assign PE_97_clock = clock;
  assign PE_97_reset = reset;
  assign PE_97_io_data_2_in_valid = PENetwork_34_io_to_pes_9_in_valid; // @[pe.scala 262:34]
  assign PE_97_io_data_2_in_bits = PENetwork_34_io_to_pes_9_in_bits; // @[pe.scala 262:34]
  assign PE_97_io_data_2_sig_stat2trans = PENetwork_34_io_to_pes_9_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_97_io_data_2_out_ready = PENetwork_34_io_to_pes_9_out_ready; // @[pe.scala 268:49]
  assign PE_97_io_data_1_in_valid = PENetwork_19_io_to_pes_9_in_valid; // @[pe.scala 262:34]
  assign PE_97_io_data_1_in_bits = PENetwork_19_io_to_pes_9_in_bits; // @[pe.scala 262:34]
  assign PE_97_io_data_0_in_valid = PENetwork_9_io_to_pes_8_in_valid; // @[pe.scala 262:34]
  assign PE_97_io_data_0_in_bits = PENetwork_9_io_to_pes_8_in_bits; // @[pe.scala 262:34]
  assign PE_98_clock = clock;
  assign PE_98_reset = reset;
  assign PE_98_io_data_2_in_valid = PENetwork_34_io_to_pes_10_in_valid; // @[pe.scala 262:34]
  assign PE_98_io_data_2_in_bits = PENetwork_34_io_to_pes_10_in_bits; // @[pe.scala 262:34]
  assign PE_98_io_data_2_sig_stat2trans = PENetwork_34_io_to_pes_10_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_98_io_data_2_out_ready = 1'h1; // @[pe.scala 268:49]
  assign PE_98_io_data_1_in_valid = PENetwork_19_io_to_pes_10_in_valid; // @[pe.scala 262:34]
  assign PE_98_io_data_1_in_bits = PENetwork_19_io_to_pes_10_in_bits; // @[pe.scala 262:34]
  assign PE_98_io_data_0_in_valid = PENetwork_10_io_to_pes_8_in_valid; // @[pe.scala 262:34]
  assign PE_98_io_data_0_in_bits = PENetwork_10_io_to_pes_8_in_bits; // @[pe.scala 262:34]
  assign PE_99_clock = clock;
  assign PE_99_reset = reset;
  assign PE_99_io_data_2_in_valid = 1'h0; // @[pe.scala 262:34]
  assign PE_99_io_data_2_in_bits = 256'h0; // @[pe.scala 262:34]
  assign PE_99_io_data_2_sig_stat2trans = PENetwork_35_io_to_pes_0_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_99_io_data_2_out_ready = PENetwork_35_io_to_pes_0_out_ready; // @[pe.scala 268:49]
  assign PE_99_io_data_1_in_valid = PENetwork_20_io_to_pes_0_in_valid; // @[pe.scala 262:34]
  assign PE_99_io_data_1_in_bits = PENetwork_20_io_to_pes_0_in_bits; // @[pe.scala 262:34]
  assign PE_99_io_data_0_in_valid = PENetwork_io_to_pes_9_in_valid; // @[pe.scala 262:34]
  assign PE_99_io_data_0_in_bits = PENetwork_io_to_pes_9_in_bits; // @[pe.scala 262:34]
  assign PE_100_clock = clock;
  assign PE_100_reset = reset;
  assign PE_100_io_data_2_in_valid = PENetwork_35_io_to_pes_1_in_valid; // @[pe.scala 262:34]
  assign PE_100_io_data_2_in_bits = PENetwork_35_io_to_pes_1_in_bits; // @[pe.scala 262:34]
  assign PE_100_io_data_2_sig_stat2trans = PENetwork_35_io_to_pes_1_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_100_io_data_2_out_ready = PENetwork_35_io_to_pes_1_out_ready; // @[pe.scala 268:49]
  assign PE_100_io_data_1_in_valid = PENetwork_20_io_to_pes_1_in_valid; // @[pe.scala 262:34]
  assign PE_100_io_data_1_in_bits = PENetwork_20_io_to_pes_1_in_bits; // @[pe.scala 262:34]
  assign PE_100_io_data_0_in_valid = PENetwork_1_io_to_pes_9_in_valid; // @[pe.scala 262:34]
  assign PE_100_io_data_0_in_bits = PENetwork_1_io_to_pes_9_in_bits; // @[pe.scala 262:34]
  assign PE_101_clock = clock;
  assign PE_101_reset = reset;
  assign PE_101_io_data_2_in_valid = PENetwork_35_io_to_pes_2_in_valid; // @[pe.scala 262:34]
  assign PE_101_io_data_2_in_bits = PENetwork_35_io_to_pes_2_in_bits; // @[pe.scala 262:34]
  assign PE_101_io_data_2_sig_stat2trans = PENetwork_35_io_to_pes_2_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_101_io_data_2_out_ready = PENetwork_35_io_to_pes_2_out_ready; // @[pe.scala 268:49]
  assign PE_101_io_data_1_in_valid = PENetwork_20_io_to_pes_2_in_valid; // @[pe.scala 262:34]
  assign PE_101_io_data_1_in_bits = PENetwork_20_io_to_pes_2_in_bits; // @[pe.scala 262:34]
  assign PE_101_io_data_0_in_valid = PENetwork_2_io_to_pes_9_in_valid; // @[pe.scala 262:34]
  assign PE_101_io_data_0_in_bits = PENetwork_2_io_to_pes_9_in_bits; // @[pe.scala 262:34]
  assign PE_102_clock = clock;
  assign PE_102_reset = reset;
  assign PE_102_io_data_2_in_valid = PENetwork_35_io_to_pes_3_in_valid; // @[pe.scala 262:34]
  assign PE_102_io_data_2_in_bits = PENetwork_35_io_to_pes_3_in_bits; // @[pe.scala 262:34]
  assign PE_102_io_data_2_sig_stat2trans = PENetwork_35_io_to_pes_3_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_102_io_data_2_out_ready = PENetwork_35_io_to_pes_3_out_ready; // @[pe.scala 268:49]
  assign PE_102_io_data_1_in_valid = PENetwork_20_io_to_pes_3_in_valid; // @[pe.scala 262:34]
  assign PE_102_io_data_1_in_bits = PENetwork_20_io_to_pes_3_in_bits; // @[pe.scala 262:34]
  assign PE_102_io_data_0_in_valid = PENetwork_3_io_to_pes_9_in_valid; // @[pe.scala 262:34]
  assign PE_102_io_data_0_in_bits = PENetwork_3_io_to_pes_9_in_bits; // @[pe.scala 262:34]
  assign PE_103_clock = clock;
  assign PE_103_reset = reset;
  assign PE_103_io_data_2_in_valid = PENetwork_35_io_to_pes_4_in_valid; // @[pe.scala 262:34]
  assign PE_103_io_data_2_in_bits = PENetwork_35_io_to_pes_4_in_bits; // @[pe.scala 262:34]
  assign PE_103_io_data_2_sig_stat2trans = PENetwork_35_io_to_pes_4_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_103_io_data_2_out_ready = PENetwork_35_io_to_pes_4_out_ready; // @[pe.scala 268:49]
  assign PE_103_io_data_1_in_valid = PENetwork_20_io_to_pes_4_in_valid; // @[pe.scala 262:34]
  assign PE_103_io_data_1_in_bits = PENetwork_20_io_to_pes_4_in_bits; // @[pe.scala 262:34]
  assign PE_103_io_data_0_in_valid = PENetwork_4_io_to_pes_9_in_valid; // @[pe.scala 262:34]
  assign PE_103_io_data_0_in_bits = PENetwork_4_io_to_pes_9_in_bits; // @[pe.scala 262:34]
  assign PE_104_clock = clock;
  assign PE_104_reset = reset;
  assign PE_104_io_data_2_in_valid = PENetwork_35_io_to_pes_5_in_valid; // @[pe.scala 262:34]
  assign PE_104_io_data_2_in_bits = PENetwork_35_io_to_pes_5_in_bits; // @[pe.scala 262:34]
  assign PE_104_io_data_2_sig_stat2trans = PENetwork_35_io_to_pes_5_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_104_io_data_2_out_ready = PENetwork_35_io_to_pes_5_out_ready; // @[pe.scala 268:49]
  assign PE_104_io_data_1_in_valid = PENetwork_20_io_to_pes_5_in_valid; // @[pe.scala 262:34]
  assign PE_104_io_data_1_in_bits = PENetwork_20_io_to_pes_5_in_bits; // @[pe.scala 262:34]
  assign PE_104_io_data_0_in_valid = PENetwork_5_io_to_pes_9_in_valid; // @[pe.scala 262:34]
  assign PE_104_io_data_0_in_bits = PENetwork_5_io_to_pes_9_in_bits; // @[pe.scala 262:34]
  assign PE_105_clock = clock;
  assign PE_105_reset = reset;
  assign PE_105_io_data_2_in_valid = PENetwork_35_io_to_pes_6_in_valid; // @[pe.scala 262:34]
  assign PE_105_io_data_2_in_bits = PENetwork_35_io_to_pes_6_in_bits; // @[pe.scala 262:34]
  assign PE_105_io_data_2_sig_stat2trans = PENetwork_35_io_to_pes_6_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_105_io_data_2_out_ready = PENetwork_35_io_to_pes_6_out_ready; // @[pe.scala 268:49]
  assign PE_105_io_data_1_in_valid = PENetwork_20_io_to_pes_6_in_valid; // @[pe.scala 262:34]
  assign PE_105_io_data_1_in_bits = PENetwork_20_io_to_pes_6_in_bits; // @[pe.scala 262:34]
  assign PE_105_io_data_0_in_valid = PENetwork_6_io_to_pes_9_in_valid; // @[pe.scala 262:34]
  assign PE_105_io_data_0_in_bits = PENetwork_6_io_to_pes_9_in_bits; // @[pe.scala 262:34]
  assign PE_106_clock = clock;
  assign PE_106_reset = reset;
  assign PE_106_io_data_2_in_valid = PENetwork_35_io_to_pes_7_in_valid; // @[pe.scala 262:34]
  assign PE_106_io_data_2_in_bits = PENetwork_35_io_to_pes_7_in_bits; // @[pe.scala 262:34]
  assign PE_106_io_data_2_sig_stat2trans = PENetwork_35_io_to_pes_7_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_106_io_data_2_out_ready = PENetwork_35_io_to_pes_7_out_ready; // @[pe.scala 268:49]
  assign PE_106_io_data_1_in_valid = PENetwork_20_io_to_pes_7_in_valid; // @[pe.scala 262:34]
  assign PE_106_io_data_1_in_bits = PENetwork_20_io_to_pes_7_in_bits; // @[pe.scala 262:34]
  assign PE_106_io_data_0_in_valid = PENetwork_7_io_to_pes_9_in_valid; // @[pe.scala 262:34]
  assign PE_106_io_data_0_in_bits = PENetwork_7_io_to_pes_9_in_bits; // @[pe.scala 262:34]
  assign PE_107_clock = clock;
  assign PE_107_reset = reset;
  assign PE_107_io_data_2_in_valid = PENetwork_35_io_to_pes_8_in_valid; // @[pe.scala 262:34]
  assign PE_107_io_data_2_in_bits = PENetwork_35_io_to_pes_8_in_bits; // @[pe.scala 262:34]
  assign PE_107_io_data_2_sig_stat2trans = PENetwork_35_io_to_pes_8_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_107_io_data_2_out_ready = PENetwork_35_io_to_pes_8_out_ready; // @[pe.scala 268:49]
  assign PE_107_io_data_1_in_valid = PENetwork_20_io_to_pes_8_in_valid; // @[pe.scala 262:34]
  assign PE_107_io_data_1_in_bits = PENetwork_20_io_to_pes_8_in_bits; // @[pe.scala 262:34]
  assign PE_107_io_data_0_in_valid = PENetwork_8_io_to_pes_9_in_valid; // @[pe.scala 262:34]
  assign PE_107_io_data_0_in_bits = PENetwork_8_io_to_pes_9_in_bits; // @[pe.scala 262:34]
  assign PE_108_clock = clock;
  assign PE_108_reset = reset;
  assign PE_108_io_data_2_in_valid = PENetwork_35_io_to_pes_9_in_valid; // @[pe.scala 262:34]
  assign PE_108_io_data_2_in_bits = PENetwork_35_io_to_pes_9_in_bits; // @[pe.scala 262:34]
  assign PE_108_io_data_2_sig_stat2trans = PENetwork_35_io_to_pes_9_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_108_io_data_2_out_ready = PENetwork_35_io_to_pes_9_out_ready; // @[pe.scala 268:49]
  assign PE_108_io_data_1_in_valid = PENetwork_20_io_to_pes_9_in_valid; // @[pe.scala 262:34]
  assign PE_108_io_data_1_in_bits = PENetwork_20_io_to_pes_9_in_bits; // @[pe.scala 262:34]
  assign PE_108_io_data_0_in_valid = PENetwork_9_io_to_pes_9_in_valid; // @[pe.scala 262:34]
  assign PE_108_io_data_0_in_bits = PENetwork_9_io_to_pes_9_in_bits; // @[pe.scala 262:34]
  assign PE_109_clock = clock;
  assign PE_109_reset = reset;
  assign PE_109_io_data_2_in_valid = PENetwork_35_io_to_pes_10_in_valid; // @[pe.scala 262:34]
  assign PE_109_io_data_2_in_bits = PENetwork_35_io_to_pes_10_in_bits; // @[pe.scala 262:34]
  assign PE_109_io_data_2_sig_stat2trans = PENetwork_35_io_to_pes_10_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_109_io_data_2_out_ready = 1'h1; // @[pe.scala 268:49]
  assign PE_109_io_data_1_in_valid = PENetwork_20_io_to_pes_10_in_valid; // @[pe.scala 262:34]
  assign PE_109_io_data_1_in_bits = PENetwork_20_io_to_pes_10_in_bits; // @[pe.scala 262:34]
  assign PE_109_io_data_0_in_valid = PENetwork_10_io_to_pes_9_in_valid; // @[pe.scala 262:34]
  assign PE_109_io_data_0_in_bits = PENetwork_10_io_to_pes_9_in_bits; // @[pe.scala 262:34]
  assign PE_110_clock = clock;
  assign PE_110_reset = reset;
  assign PE_110_io_data_2_in_valid = 1'h0; // @[pe.scala 262:34]
  assign PE_110_io_data_2_in_bits = 256'h0; // @[pe.scala 262:34]
  assign PE_110_io_data_2_sig_stat2trans = PENetwork_36_io_to_pes_0_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_110_io_data_2_out_ready = PENetwork_36_io_to_pes_0_out_ready; // @[pe.scala 268:49]
  assign PE_110_io_data_1_in_valid = PENetwork_21_io_to_pes_0_in_valid; // @[pe.scala 262:34]
  assign PE_110_io_data_1_in_bits = PENetwork_21_io_to_pes_0_in_bits; // @[pe.scala 262:34]
  assign PE_110_io_data_0_in_valid = PENetwork_io_to_pes_10_in_valid; // @[pe.scala 262:34]
  assign PE_110_io_data_0_in_bits = PENetwork_io_to_pes_10_in_bits; // @[pe.scala 262:34]
  assign PE_111_clock = clock;
  assign PE_111_reset = reset;
  assign PE_111_io_data_2_in_valid = PENetwork_36_io_to_pes_1_in_valid; // @[pe.scala 262:34]
  assign PE_111_io_data_2_in_bits = PENetwork_36_io_to_pes_1_in_bits; // @[pe.scala 262:34]
  assign PE_111_io_data_2_sig_stat2trans = PENetwork_36_io_to_pes_1_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_111_io_data_2_out_ready = PENetwork_36_io_to_pes_1_out_ready; // @[pe.scala 268:49]
  assign PE_111_io_data_1_in_valid = PENetwork_21_io_to_pes_1_in_valid; // @[pe.scala 262:34]
  assign PE_111_io_data_1_in_bits = PENetwork_21_io_to_pes_1_in_bits; // @[pe.scala 262:34]
  assign PE_111_io_data_0_in_valid = PENetwork_1_io_to_pes_10_in_valid; // @[pe.scala 262:34]
  assign PE_111_io_data_0_in_bits = PENetwork_1_io_to_pes_10_in_bits; // @[pe.scala 262:34]
  assign PE_112_clock = clock;
  assign PE_112_reset = reset;
  assign PE_112_io_data_2_in_valid = PENetwork_36_io_to_pes_2_in_valid; // @[pe.scala 262:34]
  assign PE_112_io_data_2_in_bits = PENetwork_36_io_to_pes_2_in_bits; // @[pe.scala 262:34]
  assign PE_112_io_data_2_sig_stat2trans = PENetwork_36_io_to_pes_2_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_112_io_data_2_out_ready = PENetwork_36_io_to_pes_2_out_ready; // @[pe.scala 268:49]
  assign PE_112_io_data_1_in_valid = PENetwork_21_io_to_pes_2_in_valid; // @[pe.scala 262:34]
  assign PE_112_io_data_1_in_bits = PENetwork_21_io_to_pes_2_in_bits; // @[pe.scala 262:34]
  assign PE_112_io_data_0_in_valid = PENetwork_2_io_to_pes_10_in_valid; // @[pe.scala 262:34]
  assign PE_112_io_data_0_in_bits = PENetwork_2_io_to_pes_10_in_bits; // @[pe.scala 262:34]
  assign PE_113_clock = clock;
  assign PE_113_reset = reset;
  assign PE_113_io_data_2_in_valid = PENetwork_36_io_to_pes_3_in_valid; // @[pe.scala 262:34]
  assign PE_113_io_data_2_in_bits = PENetwork_36_io_to_pes_3_in_bits; // @[pe.scala 262:34]
  assign PE_113_io_data_2_sig_stat2trans = PENetwork_36_io_to_pes_3_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_113_io_data_2_out_ready = PENetwork_36_io_to_pes_3_out_ready; // @[pe.scala 268:49]
  assign PE_113_io_data_1_in_valid = PENetwork_21_io_to_pes_3_in_valid; // @[pe.scala 262:34]
  assign PE_113_io_data_1_in_bits = PENetwork_21_io_to_pes_3_in_bits; // @[pe.scala 262:34]
  assign PE_113_io_data_0_in_valid = PENetwork_3_io_to_pes_10_in_valid; // @[pe.scala 262:34]
  assign PE_113_io_data_0_in_bits = PENetwork_3_io_to_pes_10_in_bits; // @[pe.scala 262:34]
  assign PE_114_clock = clock;
  assign PE_114_reset = reset;
  assign PE_114_io_data_2_in_valid = PENetwork_36_io_to_pes_4_in_valid; // @[pe.scala 262:34]
  assign PE_114_io_data_2_in_bits = PENetwork_36_io_to_pes_4_in_bits; // @[pe.scala 262:34]
  assign PE_114_io_data_2_sig_stat2trans = PENetwork_36_io_to_pes_4_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_114_io_data_2_out_ready = PENetwork_36_io_to_pes_4_out_ready; // @[pe.scala 268:49]
  assign PE_114_io_data_1_in_valid = PENetwork_21_io_to_pes_4_in_valid; // @[pe.scala 262:34]
  assign PE_114_io_data_1_in_bits = PENetwork_21_io_to_pes_4_in_bits; // @[pe.scala 262:34]
  assign PE_114_io_data_0_in_valid = PENetwork_4_io_to_pes_10_in_valid; // @[pe.scala 262:34]
  assign PE_114_io_data_0_in_bits = PENetwork_4_io_to_pes_10_in_bits; // @[pe.scala 262:34]
  assign PE_115_clock = clock;
  assign PE_115_reset = reset;
  assign PE_115_io_data_2_in_valid = PENetwork_36_io_to_pes_5_in_valid; // @[pe.scala 262:34]
  assign PE_115_io_data_2_in_bits = PENetwork_36_io_to_pes_5_in_bits; // @[pe.scala 262:34]
  assign PE_115_io_data_2_sig_stat2trans = PENetwork_36_io_to_pes_5_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_115_io_data_2_out_ready = PENetwork_36_io_to_pes_5_out_ready; // @[pe.scala 268:49]
  assign PE_115_io_data_1_in_valid = PENetwork_21_io_to_pes_5_in_valid; // @[pe.scala 262:34]
  assign PE_115_io_data_1_in_bits = PENetwork_21_io_to_pes_5_in_bits; // @[pe.scala 262:34]
  assign PE_115_io_data_0_in_valid = PENetwork_5_io_to_pes_10_in_valid; // @[pe.scala 262:34]
  assign PE_115_io_data_0_in_bits = PENetwork_5_io_to_pes_10_in_bits; // @[pe.scala 262:34]
  assign PE_116_clock = clock;
  assign PE_116_reset = reset;
  assign PE_116_io_data_2_in_valid = PENetwork_36_io_to_pes_6_in_valid; // @[pe.scala 262:34]
  assign PE_116_io_data_2_in_bits = PENetwork_36_io_to_pes_6_in_bits; // @[pe.scala 262:34]
  assign PE_116_io_data_2_sig_stat2trans = PENetwork_36_io_to_pes_6_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_116_io_data_2_out_ready = PENetwork_36_io_to_pes_6_out_ready; // @[pe.scala 268:49]
  assign PE_116_io_data_1_in_valid = PENetwork_21_io_to_pes_6_in_valid; // @[pe.scala 262:34]
  assign PE_116_io_data_1_in_bits = PENetwork_21_io_to_pes_6_in_bits; // @[pe.scala 262:34]
  assign PE_116_io_data_0_in_valid = PENetwork_6_io_to_pes_10_in_valid; // @[pe.scala 262:34]
  assign PE_116_io_data_0_in_bits = PENetwork_6_io_to_pes_10_in_bits; // @[pe.scala 262:34]
  assign PE_117_clock = clock;
  assign PE_117_reset = reset;
  assign PE_117_io_data_2_in_valid = PENetwork_36_io_to_pes_7_in_valid; // @[pe.scala 262:34]
  assign PE_117_io_data_2_in_bits = PENetwork_36_io_to_pes_7_in_bits; // @[pe.scala 262:34]
  assign PE_117_io_data_2_sig_stat2trans = PENetwork_36_io_to_pes_7_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_117_io_data_2_out_ready = PENetwork_36_io_to_pes_7_out_ready; // @[pe.scala 268:49]
  assign PE_117_io_data_1_in_valid = PENetwork_21_io_to_pes_7_in_valid; // @[pe.scala 262:34]
  assign PE_117_io_data_1_in_bits = PENetwork_21_io_to_pes_7_in_bits; // @[pe.scala 262:34]
  assign PE_117_io_data_0_in_valid = PENetwork_7_io_to_pes_10_in_valid; // @[pe.scala 262:34]
  assign PE_117_io_data_0_in_bits = PENetwork_7_io_to_pes_10_in_bits; // @[pe.scala 262:34]
  assign PE_118_clock = clock;
  assign PE_118_reset = reset;
  assign PE_118_io_data_2_in_valid = PENetwork_36_io_to_pes_8_in_valid; // @[pe.scala 262:34]
  assign PE_118_io_data_2_in_bits = PENetwork_36_io_to_pes_8_in_bits; // @[pe.scala 262:34]
  assign PE_118_io_data_2_sig_stat2trans = PENetwork_36_io_to_pes_8_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_118_io_data_2_out_ready = PENetwork_36_io_to_pes_8_out_ready; // @[pe.scala 268:49]
  assign PE_118_io_data_1_in_valid = PENetwork_21_io_to_pes_8_in_valid; // @[pe.scala 262:34]
  assign PE_118_io_data_1_in_bits = PENetwork_21_io_to_pes_8_in_bits; // @[pe.scala 262:34]
  assign PE_118_io_data_0_in_valid = PENetwork_8_io_to_pes_10_in_valid; // @[pe.scala 262:34]
  assign PE_118_io_data_0_in_bits = PENetwork_8_io_to_pes_10_in_bits; // @[pe.scala 262:34]
  assign PE_119_clock = clock;
  assign PE_119_reset = reset;
  assign PE_119_io_data_2_in_valid = PENetwork_36_io_to_pes_9_in_valid; // @[pe.scala 262:34]
  assign PE_119_io_data_2_in_bits = PENetwork_36_io_to_pes_9_in_bits; // @[pe.scala 262:34]
  assign PE_119_io_data_2_sig_stat2trans = PENetwork_36_io_to_pes_9_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_119_io_data_2_out_ready = PENetwork_36_io_to_pes_9_out_ready; // @[pe.scala 268:49]
  assign PE_119_io_data_1_in_valid = PENetwork_21_io_to_pes_9_in_valid; // @[pe.scala 262:34]
  assign PE_119_io_data_1_in_bits = PENetwork_21_io_to_pes_9_in_bits; // @[pe.scala 262:34]
  assign PE_119_io_data_0_in_valid = PENetwork_9_io_to_pes_10_in_valid; // @[pe.scala 262:34]
  assign PE_119_io_data_0_in_bits = PENetwork_9_io_to_pes_10_in_bits; // @[pe.scala 262:34]
  assign PE_120_clock = clock;
  assign PE_120_reset = reset;
  assign PE_120_io_data_2_in_valid = PENetwork_36_io_to_pes_10_in_valid; // @[pe.scala 262:34]
  assign PE_120_io_data_2_in_bits = PENetwork_36_io_to_pes_10_in_bits; // @[pe.scala 262:34]
  assign PE_120_io_data_2_sig_stat2trans = PENetwork_36_io_to_pes_10_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_120_io_data_2_out_ready = 1'h1; // @[pe.scala 268:49]
  assign PE_120_io_data_1_in_valid = PENetwork_21_io_to_pes_10_in_valid; // @[pe.scala 262:34]
  assign PE_120_io_data_1_in_bits = PENetwork_21_io_to_pes_10_in_bits; // @[pe.scala 262:34]
  assign PE_120_io_data_0_in_valid = PENetwork_10_io_to_pes_10_in_valid; // @[pe.scala 262:34]
  assign PE_120_io_data_0_in_bits = PENetwork_10_io_to_pes_10_in_bits; // @[pe.scala 262:34]
  assign PE_121_clock = clock;
  assign PE_121_reset = reset;
  assign PE_121_io_data_2_in_valid = 1'h0; // @[pe.scala 262:34]
  assign PE_121_io_data_2_in_bits = 256'h0; // @[pe.scala 262:34]
  assign PE_121_io_data_2_sig_stat2trans = PENetwork_37_io_to_pes_0_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_121_io_data_2_out_ready = PENetwork_37_io_to_pes_0_out_ready; // @[pe.scala 268:49]
  assign PE_121_io_data_1_in_valid = PENetwork_22_io_to_pes_0_in_valid; // @[pe.scala 262:34]
  assign PE_121_io_data_1_in_bits = PENetwork_22_io_to_pes_0_in_bits; // @[pe.scala 262:34]
  assign PE_121_io_data_0_in_valid = PENetwork_io_to_pes_11_in_valid; // @[pe.scala 262:34]
  assign PE_121_io_data_0_in_bits = PENetwork_io_to_pes_11_in_bits; // @[pe.scala 262:34]
  assign PE_122_clock = clock;
  assign PE_122_reset = reset;
  assign PE_122_io_data_2_in_valid = PENetwork_37_io_to_pes_1_in_valid; // @[pe.scala 262:34]
  assign PE_122_io_data_2_in_bits = PENetwork_37_io_to_pes_1_in_bits; // @[pe.scala 262:34]
  assign PE_122_io_data_2_sig_stat2trans = PENetwork_37_io_to_pes_1_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_122_io_data_2_out_ready = PENetwork_37_io_to_pes_1_out_ready; // @[pe.scala 268:49]
  assign PE_122_io_data_1_in_valid = PENetwork_22_io_to_pes_1_in_valid; // @[pe.scala 262:34]
  assign PE_122_io_data_1_in_bits = PENetwork_22_io_to_pes_1_in_bits; // @[pe.scala 262:34]
  assign PE_122_io_data_0_in_valid = PENetwork_1_io_to_pes_11_in_valid; // @[pe.scala 262:34]
  assign PE_122_io_data_0_in_bits = PENetwork_1_io_to_pes_11_in_bits; // @[pe.scala 262:34]
  assign PE_123_clock = clock;
  assign PE_123_reset = reset;
  assign PE_123_io_data_2_in_valid = PENetwork_37_io_to_pes_2_in_valid; // @[pe.scala 262:34]
  assign PE_123_io_data_2_in_bits = PENetwork_37_io_to_pes_2_in_bits; // @[pe.scala 262:34]
  assign PE_123_io_data_2_sig_stat2trans = PENetwork_37_io_to_pes_2_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_123_io_data_2_out_ready = PENetwork_37_io_to_pes_2_out_ready; // @[pe.scala 268:49]
  assign PE_123_io_data_1_in_valid = PENetwork_22_io_to_pes_2_in_valid; // @[pe.scala 262:34]
  assign PE_123_io_data_1_in_bits = PENetwork_22_io_to_pes_2_in_bits; // @[pe.scala 262:34]
  assign PE_123_io_data_0_in_valid = PENetwork_2_io_to_pes_11_in_valid; // @[pe.scala 262:34]
  assign PE_123_io_data_0_in_bits = PENetwork_2_io_to_pes_11_in_bits; // @[pe.scala 262:34]
  assign PE_124_clock = clock;
  assign PE_124_reset = reset;
  assign PE_124_io_data_2_in_valid = PENetwork_37_io_to_pes_3_in_valid; // @[pe.scala 262:34]
  assign PE_124_io_data_2_in_bits = PENetwork_37_io_to_pes_3_in_bits; // @[pe.scala 262:34]
  assign PE_124_io_data_2_sig_stat2trans = PENetwork_37_io_to_pes_3_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_124_io_data_2_out_ready = PENetwork_37_io_to_pes_3_out_ready; // @[pe.scala 268:49]
  assign PE_124_io_data_1_in_valid = PENetwork_22_io_to_pes_3_in_valid; // @[pe.scala 262:34]
  assign PE_124_io_data_1_in_bits = PENetwork_22_io_to_pes_3_in_bits; // @[pe.scala 262:34]
  assign PE_124_io_data_0_in_valid = PENetwork_3_io_to_pes_11_in_valid; // @[pe.scala 262:34]
  assign PE_124_io_data_0_in_bits = PENetwork_3_io_to_pes_11_in_bits; // @[pe.scala 262:34]
  assign PE_125_clock = clock;
  assign PE_125_reset = reset;
  assign PE_125_io_data_2_in_valid = PENetwork_37_io_to_pes_4_in_valid; // @[pe.scala 262:34]
  assign PE_125_io_data_2_in_bits = PENetwork_37_io_to_pes_4_in_bits; // @[pe.scala 262:34]
  assign PE_125_io_data_2_sig_stat2trans = PENetwork_37_io_to_pes_4_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_125_io_data_2_out_ready = PENetwork_37_io_to_pes_4_out_ready; // @[pe.scala 268:49]
  assign PE_125_io_data_1_in_valid = PENetwork_22_io_to_pes_4_in_valid; // @[pe.scala 262:34]
  assign PE_125_io_data_1_in_bits = PENetwork_22_io_to_pes_4_in_bits; // @[pe.scala 262:34]
  assign PE_125_io_data_0_in_valid = PENetwork_4_io_to_pes_11_in_valid; // @[pe.scala 262:34]
  assign PE_125_io_data_0_in_bits = PENetwork_4_io_to_pes_11_in_bits; // @[pe.scala 262:34]
  assign PE_126_clock = clock;
  assign PE_126_reset = reset;
  assign PE_126_io_data_2_in_valid = PENetwork_37_io_to_pes_5_in_valid; // @[pe.scala 262:34]
  assign PE_126_io_data_2_in_bits = PENetwork_37_io_to_pes_5_in_bits; // @[pe.scala 262:34]
  assign PE_126_io_data_2_sig_stat2trans = PENetwork_37_io_to_pes_5_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_126_io_data_2_out_ready = PENetwork_37_io_to_pes_5_out_ready; // @[pe.scala 268:49]
  assign PE_126_io_data_1_in_valid = PENetwork_22_io_to_pes_5_in_valid; // @[pe.scala 262:34]
  assign PE_126_io_data_1_in_bits = PENetwork_22_io_to_pes_5_in_bits; // @[pe.scala 262:34]
  assign PE_126_io_data_0_in_valid = PENetwork_5_io_to_pes_11_in_valid; // @[pe.scala 262:34]
  assign PE_126_io_data_0_in_bits = PENetwork_5_io_to_pes_11_in_bits; // @[pe.scala 262:34]
  assign PE_127_clock = clock;
  assign PE_127_reset = reset;
  assign PE_127_io_data_2_in_valid = PENetwork_37_io_to_pes_6_in_valid; // @[pe.scala 262:34]
  assign PE_127_io_data_2_in_bits = PENetwork_37_io_to_pes_6_in_bits; // @[pe.scala 262:34]
  assign PE_127_io_data_2_sig_stat2trans = PENetwork_37_io_to_pes_6_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_127_io_data_2_out_ready = PENetwork_37_io_to_pes_6_out_ready; // @[pe.scala 268:49]
  assign PE_127_io_data_1_in_valid = PENetwork_22_io_to_pes_6_in_valid; // @[pe.scala 262:34]
  assign PE_127_io_data_1_in_bits = PENetwork_22_io_to_pes_6_in_bits; // @[pe.scala 262:34]
  assign PE_127_io_data_0_in_valid = PENetwork_6_io_to_pes_11_in_valid; // @[pe.scala 262:34]
  assign PE_127_io_data_0_in_bits = PENetwork_6_io_to_pes_11_in_bits; // @[pe.scala 262:34]
  assign PE_128_clock = clock;
  assign PE_128_reset = reset;
  assign PE_128_io_data_2_in_valid = PENetwork_37_io_to_pes_7_in_valid; // @[pe.scala 262:34]
  assign PE_128_io_data_2_in_bits = PENetwork_37_io_to_pes_7_in_bits; // @[pe.scala 262:34]
  assign PE_128_io_data_2_sig_stat2trans = PENetwork_37_io_to_pes_7_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_128_io_data_2_out_ready = PENetwork_37_io_to_pes_7_out_ready; // @[pe.scala 268:49]
  assign PE_128_io_data_1_in_valid = PENetwork_22_io_to_pes_7_in_valid; // @[pe.scala 262:34]
  assign PE_128_io_data_1_in_bits = PENetwork_22_io_to_pes_7_in_bits; // @[pe.scala 262:34]
  assign PE_128_io_data_0_in_valid = PENetwork_7_io_to_pes_11_in_valid; // @[pe.scala 262:34]
  assign PE_128_io_data_0_in_bits = PENetwork_7_io_to_pes_11_in_bits; // @[pe.scala 262:34]
  assign PE_129_clock = clock;
  assign PE_129_reset = reset;
  assign PE_129_io_data_2_in_valid = PENetwork_37_io_to_pes_8_in_valid; // @[pe.scala 262:34]
  assign PE_129_io_data_2_in_bits = PENetwork_37_io_to_pes_8_in_bits; // @[pe.scala 262:34]
  assign PE_129_io_data_2_sig_stat2trans = PENetwork_37_io_to_pes_8_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_129_io_data_2_out_ready = PENetwork_37_io_to_pes_8_out_ready; // @[pe.scala 268:49]
  assign PE_129_io_data_1_in_valid = PENetwork_22_io_to_pes_8_in_valid; // @[pe.scala 262:34]
  assign PE_129_io_data_1_in_bits = PENetwork_22_io_to_pes_8_in_bits; // @[pe.scala 262:34]
  assign PE_129_io_data_0_in_valid = PENetwork_8_io_to_pes_11_in_valid; // @[pe.scala 262:34]
  assign PE_129_io_data_0_in_bits = PENetwork_8_io_to_pes_11_in_bits; // @[pe.scala 262:34]
  assign PE_130_clock = clock;
  assign PE_130_reset = reset;
  assign PE_130_io_data_2_in_valid = PENetwork_37_io_to_pes_9_in_valid; // @[pe.scala 262:34]
  assign PE_130_io_data_2_in_bits = PENetwork_37_io_to_pes_9_in_bits; // @[pe.scala 262:34]
  assign PE_130_io_data_2_sig_stat2trans = PENetwork_37_io_to_pes_9_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_130_io_data_2_out_ready = PENetwork_37_io_to_pes_9_out_ready; // @[pe.scala 268:49]
  assign PE_130_io_data_1_in_valid = PENetwork_22_io_to_pes_9_in_valid; // @[pe.scala 262:34]
  assign PE_130_io_data_1_in_bits = PENetwork_22_io_to_pes_9_in_bits; // @[pe.scala 262:34]
  assign PE_130_io_data_0_in_valid = PENetwork_9_io_to_pes_11_in_valid; // @[pe.scala 262:34]
  assign PE_130_io_data_0_in_bits = PENetwork_9_io_to_pes_11_in_bits; // @[pe.scala 262:34]
  assign PE_131_clock = clock;
  assign PE_131_reset = reset;
  assign PE_131_io_data_2_in_valid = PENetwork_37_io_to_pes_10_in_valid; // @[pe.scala 262:34]
  assign PE_131_io_data_2_in_bits = PENetwork_37_io_to_pes_10_in_bits; // @[pe.scala 262:34]
  assign PE_131_io_data_2_sig_stat2trans = PENetwork_37_io_to_pes_10_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_131_io_data_2_out_ready = 1'h1; // @[pe.scala 268:49]
  assign PE_131_io_data_1_in_valid = PENetwork_22_io_to_pes_10_in_valid; // @[pe.scala 262:34]
  assign PE_131_io_data_1_in_bits = PENetwork_22_io_to_pes_10_in_bits; // @[pe.scala 262:34]
  assign PE_131_io_data_0_in_valid = PENetwork_10_io_to_pes_11_in_valid; // @[pe.scala 262:34]
  assign PE_131_io_data_0_in_bits = PENetwork_10_io_to_pes_11_in_bits; // @[pe.scala 262:34]
  assign PE_132_clock = clock;
  assign PE_132_reset = reset;
  assign PE_132_io_data_2_in_valid = 1'h0; // @[pe.scala 262:34]
  assign PE_132_io_data_2_in_bits = 256'h0; // @[pe.scala 262:34]
  assign PE_132_io_data_2_sig_stat2trans = PENetwork_38_io_to_pes_0_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_132_io_data_2_out_ready = PENetwork_38_io_to_pes_0_out_ready; // @[pe.scala 268:49]
  assign PE_132_io_data_1_in_valid = PENetwork_23_io_to_pes_0_in_valid; // @[pe.scala 262:34]
  assign PE_132_io_data_1_in_bits = PENetwork_23_io_to_pes_0_in_bits; // @[pe.scala 262:34]
  assign PE_132_io_data_0_in_valid = PENetwork_io_to_pes_12_in_valid; // @[pe.scala 262:34]
  assign PE_132_io_data_0_in_bits = PENetwork_io_to_pes_12_in_bits; // @[pe.scala 262:34]
  assign PE_133_clock = clock;
  assign PE_133_reset = reset;
  assign PE_133_io_data_2_in_valid = PENetwork_38_io_to_pes_1_in_valid; // @[pe.scala 262:34]
  assign PE_133_io_data_2_in_bits = PENetwork_38_io_to_pes_1_in_bits; // @[pe.scala 262:34]
  assign PE_133_io_data_2_sig_stat2trans = PENetwork_38_io_to_pes_1_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_133_io_data_2_out_ready = PENetwork_38_io_to_pes_1_out_ready; // @[pe.scala 268:49]
  assign PE_133_io_data_1_in_valid = PENetwork_23_io_to_pes_1_in_valid; // @[pe.scala 262:34]
  assign PE_133_io_data_1_in_bits = PENetwork_23_io_to_pes_1_in_bits; // @[pe.scala 262:34]
  assign PE_133_io_data_0_in_valid = PENetwork_1_io_to_pes_12_in_valid; // @[pe.scala 262:34]
  assign PE_133_io_data_0_in_bits = PENetwork_1_io_to_pes_12_in_bits; // @[pe.scala 262:34]
  assign PE_134_clock = clock;
  assign PE_134_reset = reset;
  assign PE_134_io_data_2_in_valid = PENetwork_38_io_to_pes_2_in_valid; // @[pe.scala 262:34]
  assign PE_134_io_data_2_in_bits = PENetwork_38_io_to_pes_2_in_bits; // @[pe.scala 262:34]
  assign PE_134_io_data_2_sig_stat2trans = PENetwork_38_io_to_pes_2_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_134_io_data_2_out_ready = PENetwork_38_io_to_pes_2_out_ready; // @[pe.scala 268:49]
  assign PE_134_io_data_1_in_valid = PENetwork_23_io_to_pes_2_in_valid; // @[pe.scala 262:34]
  assign PE_134_io_data_1_in_bits = PENetwork_23_io_to_pes_2_in_bits; // @[pe.scala 262:34]
  assign PE_134_io_data_0_in_valid = PENetwork_2_io_to_pes_12_in_valid; // @[pe.scala 262:34]
  assign PE_134_io_data_0_in_bits = PENetwork_2_io_to_pes_12_in_bits; // @[pe.scala 262:34]
  assign PE_135_clock = clock;
  assign PE_135_reset = reset;
  assign PE_135_io_data_2_in_valid = PENetwork_38_io_to_pes_3_in_valid; // @[pe.scala 262:34]
  assign PE_135_io_data_2_in_bits = PENetwork_38_io_to_pes_3_in_bits; // @[pe.scala 262:34]
  assign PE_135_io_data_2_sig_stat2trans = PENetwork_38_io_to_pes_3_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_135_io_data_2_out_ready = PENetwork_38_io_to_pes_3_out_ready; // @[pe.scala 268:49]
  assign PE_135_io_data_1_in_valid = PENetwork_23_io_to_pes_3_in_valid; // @[pe.scala 262:34]
  assign PE_135_io_data_1_in_bits = PENetwork_23_io_to_pes_3_in_bits; // @[pe.scala 262:34]
  assign PE_135_io_data_0_in_valid = PENetwork_3_io_to_pes_12_in_valid; // @[pe.scala 262:34]
  assign PE_135_io_data_0_in_bits = PENetwork_3_io_to_pes_12_in_bits; // @[pe.scala 262:34]
  assign PE_136_clock = clock;
  assign PE_136_reset = reset;
  assign PE_136_io_data_2_in_valid = PENetwork_38_io_to_pes_4_in_valid; // @[pe.scala 262:34]
  assign PE_136_io_data_2_in_bits = PENetwork_38_io_to_pes_4_in_bits; // @[pe.scala 262:34]
  assign PE_136_io_data_2_sig_stat2trans = PENetwork_38_io_to_pes_4_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_136_io_data_2_out_ready = PENetwork_38_io_to_pes_4_out_ready; // @[pe.scala 268:49]
  assign PE_136_io_data_1_in_valid = PENetwork_23_io_to_pes_4_in_valid; // @[pe.scala 262:34]
  assign PE_136_io_data_1_in_bits = PENetwork_23_io_to_pes_4_in_bits; // @[pe.scala 262:34]
  assign PE_136_io_data_0_in_valid = PENetwork_4_io_to_pes_12_in_valid; // @[pe.scala 262:34]
  assign PE_136_io_data_0_in_bits = PENetwork_4_io_to_pes_12_in_bits; // @[pe.scala 262:34]
  assign PE_137_clock = clock;
  assign PE_137_reset = reset;
  assign PE_137_io_data_2_in_valid = PENetwork_38_io_to_pes_5_in_valid; // @[pe.scala 262:34]
  assign PE_137_io_data_2_in_bits = PENetwork_38_io_to_pes_5_in_bits; // @[pe.scala 262:34]
  assign PE_137_io_data_2_sig_stat2trans = PENetwork_38_io_to_pes_5_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_137_io_data_2_out_ready = PENetwork_38_io_to_pes_5_out_ready; // @[pe.scala 268:49]
  assign PE_137_io_data_1_in_valid = PENetwork_23_io_to_pes_5_in_valid; // @[pe.scala 262:34]
  assign PE_137_io_data_1_in_bits = PENetwork_23_io_to_pes_5_in_bits; // @[pe.scala 262:34]
  assign PE_137_io_data_0_in_valid = PENetwork_5_io_to_pes_12_in_valid; // @[pe.scala 262:34]
  assign PE_137_io_data_0_in_bits = PENetwork_5_io_to_pes_12_in_bits; // @[pe.scala 262:34]
  assign PE_138_clock = clock;
  assign PE_138_reset = reset;
  assign PE_138_io_data_2_in_valid = PENetwork_38_io_to_pes_6_in_valid; // @[pe.scala 262:34]
  assign PE_138_io_data_2_in_bits = PENetwork_38_io_to_pes_6_in_bits; // @[pe.scala 262:34]
  assign PE_138_io_data_2_sig_stat2trans = PENetwork_38_io_to_pes_6_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_138_io_data_2_out_ready = PENetwork_38_io_to_pes_6_out_ready; // @[pe.scala 268:49]
  assign PE_138_io_data_1_in_valid = PENetwork_23_io_to_pes_6_in_valid; // @[pe.scala 262:34]
  assign PE_138_io_data_1_in_bits = PENetwork_23_io_to_pes_6_in_bits; // @[pe.scala 262:34]
  assign PE_138_io_data_0_in_valid = PENetwork_6_io_to_pes_12_in_valid; // @[pe.scala 262:34]
  assign PE_138_io_data_0_in_bits = PENetwork_6_io_to_pes_12_in_bits; // @[pe.scala 262:34]
  assign PE_139_clock = clock;
  assign PE_139_reset = reset;
  assign PE_139_io_data_2_in_valid = PENetwork_38_io_to_pes_7_in_valid; // @[pe.scala 262:34]
  assign PE_139_io_data_2_in_bits = PENetwork_38_io_to_pes_7_in_bits; // @[pe.scala 262:34]
  assign PE_139_io_data_2_sig_stat2trans = PENetwork_38_io_to_pes_7_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_139_io_data_2_out_ready = PENetwork_38_io_to_pes_7_out_ready; // @[pe.scala 268:49]
  assign PE_139_io_data_1_in_valid = PENetwork_23_io_to_pes_7_in_valid; // @[pe.scala 262:34]
  assign PE_139_io_data_1_in_bits = PENetwork_23_io_to_pes_7_in_bits; // @[pe.scala 262:34]
  assign PE_139_io_data_0_in_valid = PENetwork_7_io_to_pes_12_in_valid; // @[pe.scala 262:34]
  assign PE_139_io_data_0_in_bits = PENetwork_7_io_to_pes_12_in_bits; // @[pe.scala 262:34]
  assign PE_140_clock = clock;
  assign PE_140_reset = reset;
  assign PE_140_io_data_2_in_valid = PENetwork_38_io_to_pes_8_in_valid; // @[pe.scala 262:34]
  assign PE_140_io_data_2_in_bits = PENetwork_38_io_to_pes_8_in_bits; // @[pe.scala 262:34]
  assign PE_140_io_data_2_sig_stat2trans = PENetwork_38_io_to_pes_8_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_140_io_data_2_out_ready = PENetwork_38_io_to_pes_8_out_ready; // @[pe.scala 268:49]
  assign PE_140_io_data_1_in_valid = PENetwork_23_io_to_pes_8_in_valid; // @[pe.scala 262:34]
  assign PE_140_io_data_1_in_bits = PENetwork_23_io_to_pes_8_in_bits; // @[pe.scala 262:34]
  assign PE_140_io_data_0_in_valid = PENetwork_8_io_to_pes_12_in_valid; // @[pe.scala 262:34]
  assign PE_140_io_data_0_in_bits = PENetwork_8_io_to_pes_12_in_bits; // @[pe.scala 262:34]
  assign PE_141_clock = clock;
  assign PE_141_reset = reset;
  assign PE_141_io_data_2_in_valid = PENetwork_38_io_to_pes_9_in_valid; // @[pe.scala 262:34]
  assign PE_141_io_data_2_in_bits = PENetwork_38_io_to_pes_9_in_bits; // @[pe.scala 262:34]
  assign PE_141_io_data_2_sig_stat2trans = PENetwork_38_io_to_pes_9_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_141_io_data_2_out_ready = PENetwork_38_io_to_pes_9_out_ready; // @[pe.scala 268:49]
  assign PE_141_io_data_1_in_valid = PENetwork_23_io_to_pes_9_in_valid; // @[pe.scala 262:34]
  assign PE_141_io_data_1_in_bits = PENetwork_23_io_to_pes_9_in_bits; // @[pe.scala 262:34]
  assign PE_141_io_data_0_in_valid = PENetwork_9_io_to_pes_12_in_valid; // @[pe.scala 262:34]
  assign PE_141_io_data_0_in_bits = PENetwork_9_io_to_pes_12_in_bits; // @[pe.scala 262:34]
  assign PE_142_clock = clock;
  assign PE_142_reset = reset;
  assign PE_142_io_data_2_in_valid = PENetwork_38_io_to_pes_10_in_valid; // @[pe.scala 262:34]
  assign PE_142_io_data_2_in_bits = PENetwork_38_io_to_pes_10_in_bits; // @[pe.scala 262:34]
  assign PE_142_io_data_2_sig_stat2trans = PENetwork_38_io_to_pes_10_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_142_io_data_2_out_ready = 1'h1; // @[pe.scala 268:49]
  assign PE_142_io_data_1_in_valid = PENetwork_23_io_to_pes_10_in_valid; // @[pe.scala 262:34]
  assign PE_142_io_data_1_in_bits = PENetwork_23_io_to_pes_10_in_bits; // @[pe.scala 262:34]
  assign PE_142_io_data_0_in_valid = PENetwork_10_io_to_pes_12_in_valid; // @[pe.scala 262:34]
  assign PE_142_io_data_0_in_bits = PENetwork_10_io_to_pes_12_in_bits; // @[pe.scala 262:34]
  assign PE_143_clock = clock;
  assign PE_143_reset = reset;
  assign PE_143_io_data_2_in_valid = 1'h0; // @[pe.scala 262:34]
  assign PE_143_io_data_2_in_bits = 256'h0; // @[pe.scala 262:34]
  assign PE_143_io_data_2_sig_stat2trans = PENetwork_39_io_to_pes_0_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_143_io_data_2_out_ready = PENetwork_39_io_to_pes_0_out_ready; // @[pe.scala 268:49]
  assign PE_143_io_data_1_in_valid = PENetwork_24_io_to_pes_0_in_valid; // @[pe.scala 262:34]
  assign PE_143_io_data_1_in_bits = PENetwork_24_io_to_pes_0_in_bits; // @[pe.scala 262:34]
  assign PE_143_io_data_0_in_valid = PENetwork_io_to_pes_13_in_valid; // @[pe.scala 262:34]
  assign PE_143_io_data_0_in_bits = PENetwork_io_to_pes_13_in_bits; // @[pe.scala 262:34]
  assign PE_144_clock = clock;
  assign PE_144_reset = reset;
  assign PE_144_io_data_2_in_valid = PENetwork_39_io_to_pes_1_in_valid; // @[pe.scala 262:34]
  assign PE_144_io_data_2_in_bits = PENetwork_39_io_to_pes_1_in_bits; // @[pe.scala 262:34]
  assign PE_144_io_data_2_sig_stat2trans = PENetwork_39_io_to_pes_1_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_144_io_data_2_out_ready = PENetwork_39_io_to_pes_1_out_ready; // @[pe.scala 268:49]
  assign PE_144_io_data_1_in_valid = PENetwork_24_io_to_pes_1_in_valid; // @[pe.scala 262:34]
  assign PE_144_io_data_1_in_bits = PENetwork_24_io_to_pes_1_in_bits; // @[pe.scala 262:34]
  assign PE_144_io_data_0_in_valid = PENetwork_1_io_to_pes_13_in_valid; // @[pe.scala 262:34]
  assign PE_144_io_data_0_in_bits = PENetwork_1_io_to_pes_13_in_bits; // @[pe.scala 262:34]
  assign PE_145_clock = clock;
  assign PE_145_reset = reset;
  assign PE_145_io_data_2_in_valid = PENetwork_39_io_to_pes_2_in_valid; // @[pe.scala 262:34]
  assign PE_145_io_data_2_in_bits = PENetwork_39_io_to_pes_2_in_bits; // @[pe.scala 262:34]
  assign PE_145_io_data_2_sig_stat2trans = PENetwork_39_io_to_pes_2_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_145_io_data_2_out_ready = PENetwork_39_io_to_pes_2_out_ready; // @[pe.scala 268:49]
  assign PE_145_io_data_1_in_valid = PENetwork_24_io_to_pes_2_in_valid; // @[pe.scala 262:34]
  assign PE_145_io_data_1_in_bits = PENetwork_24_io_to_pes_2_in_bits; // @[pe.scala 262:34]
  assign PE_145_io_data_0_in_valid = PENetwork_2_io_to_pes_13_in_valid; // @[pe.scala 262:34]
  assign PE_145_io_data_0_in_bits = PENetwork_2_io_to_pes_13_in_bits; // @[pe.scala 262:34]
  assign PE_146_clock = clock;
  assign PE_146_reset = reset;
  assign PE_146_io_data_2_in_valid = PENetwork_39_io_to_pes_3_in_valid; // @[pe.scala 262:34]
  assign PE_146_io_data_2_in_bits = PENetwork_39_io_to_pes_3_in_bits; // @[pe.scala 262:34]
  assign PE_146_io_data_2_sig_stat2trans = PENetwork_39_io_to_pes_3_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_146_io_data_2_out_ready = PENetwork_39_io_to_pes_3_out_ready; // @[pe.scala 268:49]
  assign PE_146_io_data_1_in_valid = PENetwork_24_io_to_pes_3_in_valid; // @[pe.scala 262:34]
  assign PE_146_io_data_1_in_bits = PENetwork_24_io_to_pes_3_in_bits; // @[pe.scala 262:34]
  assign PE_146_io_data_0_in_valid = PENetwork_3_io_to_pes_13_in_valid; // @[pe.scala 262:34]
  assign PE_146_io_data_0_in_bits = PENetwork_3_io_to_pes_13_in_bits; // @[pe.scala 262:34]
  assign PE_147_clock = clock;
  assign PE_147_reset = reset;
  assign PE_147_io_data_2_in_valid = PENetwork_39_io_to_pes_4_in_valid; // @[pe.scala 262:34]
  assign PE_147_io_data_2_in_bits = PENetwork_39_io_to_pes_4_in_bits; // @[pe.scala 262:34]
  assign PE_147_io_data_2_sig_stat2trans = PENetwork_39_io_to_pes_4_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_147_io_data_2_out_ready = PENetwork_39_io_to_pes_4_out_ready; // @[pe.scala 268:49]
  assign PE_147_io_data_1_in_valid = PENetwork_24_io_to_pes_4_in_valid; // @[pe.scala 262:34]
  assign PE_147_io_data_1_in_bits = PENetwork_24_io_to_pes_4_in_bits; // @[pe.scala 262:34]
  assign PE_147_io_data_0_in_valid = PENetwork_4_io_to_pes_13_in_valid; // @[pe.scala 262:34]
  assign PE_147_io_data_0_in_bits = PENetwork_4_io_to_pes_13_in_bits; // @[pe.scala 262:34]
  assign PE_148_clock = clock;
  assign PE_148_reset = reset;
  assign PE_148_io_data_2_in_valid = PENetwork_39_io_to_pes_5_in_valid; // @[pe.scala 262:34]
  assign PE_148_io_data_2_in_bits = PENetwork_39_io_to_pes_5_in_bits; // @[pe.scala 262:34]
  assign PE_148_io_data_2_sig_stat2trans = PENetwork_39_io_to_pes_5_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_148_io_data_2_out_ready = PENetwork_39_io_to_pes_5_out_ready; // @[pe.scala 268:49]
  assign PE_148_io_data_1_in_valid = PENetwork_24_io_to_pes_5_in_valid; // @[pe.scala 262:34]
  assign PE_148_io_data_1_in_bits = PENetwork_24_io_to_pes_5_in_bits; // @[pe.scala 262:34]
  assign PE_148_io_data_0_in_valid = PENetwork_5_io_to_pes_13_in_valid; // @[pe.scala 262:34]
  assign PE_148_io_data_0_in_bits = PENetwork_5_io_to_pes_13_in_bits; // @[pe.scala 262:34]
  assign PE_149_clock = clock;
  assign PE_149_reset = reset;
  assign PE_149_io_data_2_in_valid = PENetwork_39_io_to_pes_6_in_valid; // @[pe.scala 262:34]
  assign PE_149_io_data_2_in_bits = PENetwork_39_io_to_pes_6_in_bits; // @[pe.scala 262:34]
  assign PE_149_io_data_2_sig_stat2trans = PENetwork_39_io_to_pes_6_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_149_io_data_2_out_ready = PENetwork_39_io_to_pes_6_out_ready; // @[pe.scala 268:49]
  assign PE_149_io_data_1_in_valid = PENetwork_24_io_to_pes_6_in_valid; // @[pe.scala 262:34]
  assign PE_149_io_data_1_in_bits = PENetwork_24_io_to_pes_6_in_bits; // @[pe.scala 262:34]
  assign PE_149_io_data_0_in_valid = PENetwork_6_io_to_pes_13_in_valid; // @[pe.scala 262:34]
  assign PE_149_io_data_0_in_bits = PENetwork_6_io_to_pes_13_in_bits; // @[pe.scala 262:34]
  assign PE_150_clock = clock;
  assign PE_150_reset = reset;
  assign PE_150_io_data_2_in_valid = PENetwork_39_io_to_pes_7_in_valid; // @[pe.scala 262:34]
  assign PE_150_io_data_2_in_bits = PENetwork_39_io_to_pes_7_in_bits; // @[pe.scala 262:34]
  assign PE_150_io_data_2_sig_stat2trans = PENetwork_39_io_to_pes_7_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_150_io_data_2_out_ready = PENetwork_39_io_to_pes_7_out_ready; // @[pe.scala 268:49]
  assign PE_150_io_data_1_in_valid = PENetwork_24_io_to_pes_7_in_valid; // @[pe.scala 262:34]
  assign PE_150_io_data_1_in_bits = PENetwork_24_io_to_pes_7_in_bits; // @[pe.scala 262:34]
  assign PE_150_io_data_0_in_valid = PENetwork_7_io_to_pes_13_in_valid; // @[pe.scala 262:34]
  assign PE_150_io_data_0_in_bits = PENetwork_7_io_to_pes_13_in_bits; // @[pe.scala 262:34]
  assign PE_151_clock = clock;
  assign PE_151_reset = reset;
  assign PE_151_io_data_2_in_valid = PENetwork_39_io_to_pes_8_in_valid; // @[pe.scala 262:34]
  assign PE_151_io_data_2_in_bits = PENetwork_39_io_to_pes_8_in_bits; // @[pe.scala 262:34]
  assign PE_151_io_data_2_sig_stat2trans = PENetwork_39_io_to_pes_8_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_151_io_data_2_out_ready = PENetwork_39_io_to_pes_8_out_ready; // @[pe.scala 268:49]
  assign PE_151_io_data_1_in_valid = PENetwork_24_io_to_pes_8_in_valid; // @[pe.scala 262:34]
  assign PE_151_io_data_1_in_bits = PENetwork_24_io_to_pes_8_in_bits; // @[pe.scala 262:34]
  assign PE_151_io_data_0_in_valid = PENetwork_8_io_to_pes_13_in_valid; // @[pe.scala 262:34]
  assign PE_151_io_data_0_in_bits = PENetwork_8_io_to_pes_13_in_bits; // @[pe.scala 262:34]
  assign PE_152_clock = clock;
  assign PE_152_reset = reset;
  assign PE_152_io_data_2_in_valid = PENetwork_39_io_to_pes_9_in_valid; // @[pe.scala 262:34]
  assign PE_152_io_data_2_in_bits = PENetwork_39_io_to_pes_9_in_bits; // @[pe.scala 262:34]
  assign PE_152_io_data_2_sig_stat2trans = PENetwork_39_io_to_pes_9_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_152_io_data_2_out_ready = PENetwork_39_io_to_pes_9_out_ready; // @[pe.scala 268:49]
  assign PE_152_io_data_1_in_valid = PENetwork_24_io_to_pes_9_in_valid; // @[pe.scala 262:34]
  assign PE_152_io_data_1_in_bits = PENetwork_24_io_to_pes_9_in_bits; // @[pe.scala 262:34]
  assign PE_152_io_data_0_in_valid = PENetwork_9_io_to_pes_13_in_valid; // @[pe.scala 262:34]
  assign PE_152_io_data_0_in_bits = PENetwork_9_io_to_pes_13_in_bits; // @[pe.scala 262:34]
  assign PE_153_clock = clock;
  assign PE_153_reset = reset;
  assign PE_153_io_data_2_in_valid = PENetwork_39_io_to_pes_10_in_valid; // @[pe.scala 262:34]
  assign PE_153_io_data_2_in_bits = PENetwork_39_io_to_pes_10_in_bits; // @[pe.scala 262:34]
  assign PE_153_io_data_2_sig_stat2trans = PENetwork_39_io_to_pes_10_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_153_io_data_2_out_ready = 1'h1; // @[pe.scala 268:49]
  assign PE_153_io_data_1_in_valid = PENetwork_24_io_to_pes_10_in_valid; // @[pe.scala 262:34]
  assign PE_153_io_data_1_in_bits = PENetwork_24_io_to_pes_10_in_bits; // @[pe.scala 262:34]
  assign PE_153_io_data_0_in_valid = PENetwork_10_io_to_pes_13_in_valid; // @[pe.scala 262:34]
  assign PE_153_io_data_0_in_bits = PENetwork_10_io_to_pes_13_in_bits; // @[pe.scala 262:34]
  assign PE_154_clock = clock;
  assign PE_154_reset = reset;
  assign PE_154_io_data_2_in_valid = 1'h0; // @[pe.scala 262:34]
  assign PE_154_io_data_2_in_bits = 256'h0; // @[pe.scala 262:34]
  assign PE_154_io_data_2_sig_stat2trans = PENetwork_40_io_to_pes_0_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_154_io_data_2_out_ready = PENetwork_40_io_to_pes_0_out_ready; // @[pe.scala 268:49]
  assign PE_154_io_data_1_in_valid = PENetwork_25_io_to_pes_0_in_valid; // @[pe.scala 262:34]
  assign PE_154_io_data_1_in_bits = PENetwork_25_io_to_pes_0_in_bits; // @[pe.scala 262:34]
  assign PE_154_io_data_0_in_valid = PENetwork_io_to_pes_14_in_valid; // @[pe.scala 262:34]
  assign PE_154_io_data_0_in_bits = PENetwork_io_to_pes_14_in_bits; // @[pe.scala 262:34]
  assign PE_155_clock = clock;
  assign PE_155_reset = reset;
  assign PE_155_io_data_2_in_valid = PENetwork_40_io_to_pes_1_in_valid; // @[pe.scala 262:34]
  assign PE_155_io_data_2_in_bits = PENetwork_40_io_to_pes_1_in_bits; // @[pe.scala 262:34]
  assign PE_155_io_data_2_sig_stat2trans = PENetwork_40_io_to_pes_1_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_155_io_data_2_out_ready = PENetwork_40_io_to_pes_1_out_ready; // @[pe.scala 268:49]
  assign PE_155_io_data_1_in_valid = PENetwork_25_io_to_pes_1_in_valid; // @[pe.scala 262:34]
  assign PE_155_io_data_1_in_bits = PENetwork_25_io_to_pes_1_in_bits; // @[pe.scala 262:34]
  assign PE_155_io_data_0_in_valid = PENetwork_1_io_to_pes_14_in_valid; // @[pe.scala 262:34]
  assign PE_155_io_data_0_in_bits = PENetwork_1_io_to_pes_14_in_bits; // @[pe.scala 262:34]
  assign PE_156_clock = clock;
  assign PE_156_reset = reset;
  assign PE_156_io_data_2_in_valid = PENetwork_40_io_to_pes_2_in_valid; // @[pe.scala 262:34]
  assign PE_156_io_data_2_in_bits = PENetwork_40_io_to_pes_2_in_bits; // @[pe.scala 262:34]
  assign PE_156_io_data_2_sig_stat2trans = PENetwork_40_io_to_pes_2_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_156_io_data_2_out_ready = PENetwork_40_io_to_pes_2_out_ready; // @[pe.scala 268:49]
  assign PE_156_io_data_1_in_valid = PENetwork_25_io_to_pes_2_in_valid; // @[pe.scala 262:34]
  assign PE_156_io_data_1_in_bits = PENetwork_25_io_to_pes_2_in_bits; // @[pe.scala 262:34]
  assign PE_156_io_data_0_in_valid = PENetwork_2_io_to_pes_14_in_valid; // @[pe.scala 262:34]
  assign PE_156_io_data_0_in_bits = PENetwork_2_io_to_pes_14_in_bits; // @[pe.scala 262:34]
  assign PE_157_clock = clock;
  assign PE_157_reset = reset;
  assign PE_157_io_data_2_in_valid = PENetwork_40_io_to_pes_3_in_valid; // @[pe.scala 262:34]
  assign PE_157_io_data_2_in_bits = PENetwork_40_io_to_pes_3_in_bits; // @[pe.scala 262:34]
  assign PE_157_io_data_2_sig_stat2trans = PENetwork_40_io_to_pes_3_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_157_io_data_2_out_ready = PENetwork_40_io_to_pes_3_out_ready; // @[pe.scala 268:49]
  assign PE_157_io_data_1_in_valid = PENetwork_25_io_to_pes_3_in_valid; // @[pe.scala 262:34]
  assign PE_157_io_data_1_in_bits = PENetwork_25_io_to_pes_3_in_bits; // @[pe.scala 262:34]
  assign PE_157_io_data_0_in_valid = PENetwork_3_io_to_pes_14_in_valid; // @[pe.scala 262:34]
  assign PE_157_io_data_0_in_bits = PENetwork_3_io_to_pes_14_in_bits; // @[pe.scala 262:34]
  assign PE_158_clock = clock;
  assign PE_158_reset = reset;
  assign PE_158_io_data_2_in_valid = PENetwork_40_io_to_pes_4_in_valid; // @[pe.scala 262:34]
  assign PE_158_io_data_2_in_bits = PENetwork_40_io_to_pes_4_in_bits; // @[pe.scala 262:34]
  assign PE_158_io_data_2_sig_stat2trans = PENetwork_40_io_to_pes_4_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_158_io_data_2_out_ready = PENetwork_40_io_to_pes_4_out_ready; // @[pe.scala 268:49]
  assign PE_158_io_data_1_in_valid = PENetwork_25_io_to_pes_4_in_valid; // @[pe.scala 262:34]
  assign PE_158_io_data_1_in_bits = PENetwork_25_io_to_pes_4_in_bits; // @[pe.scala 262:34]
  assign PE_158_io_data_0_in_valid = PENetwork_4_io_to_pes_14_in_valid; // @[pe.scala 262:34]
  assign PE_158_io_data_0_in_bits = PENetwork_4_io_to_pes_14_in_bits; // @[pe.scala 262:34]
  assign PE_159_clock = clock;
  assign PE_159_reset = reset;
  assign PE_159_io_data_2_in_valid = PENetwork_40_io_to_pes_5_in_valid; // @[pe.scala 262:34]
  assign PE_159_io_data_2_in_bits = PENetwork_40_io_to_pes_5_in_bits; // @[pe.scala 262:34]
  assign PE_159_io_data_2_sig_stat2trans = PENetwork_40_io_to_pes_5_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_159_io_data_2_out_ready = PENetwork_40_io_to_pes_5_out_ready; // @[pe.scala 268:49]
  assign PE_159_io_data_1_in_valid = PENetwork_25_io_to_pes_5_in_valid; // @[pe.scala 262:34]
  assign PE_159_io_data_1_in_bits = PENetwork_25_io_to_pes_5_in_bits; // @[pe.scala 262:34]
  assign PE_159_io_data_0_in_valid = PENetwork_5_io_to_pes_14_in_valid; // @[pe.scala 262:34]
  assign PE_159_io_data_0_in_bits = PENetwork_5_io_to_pes_14_in_bits; // @[pe.scala 262:34]
  assign PE_160_clock = clock;
  assign PE_160_reset = reset;
  assign PE_160_io_data_2_in_valid = PENetwork_40_io_to_pes_6_in_valid; // @[pe.scala 262:34]
  assign PE_160_io_data_2_in_bits = PENetwork_40_io_to_pes_6_in_bits; // @[pe.scala 262:34]
  assign PE_160_io_data_2_sig_stat2trans = PENetwork_40_io_to_pes_6_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_160_io_data_2_out_ready = PENetwork_40_io_to_pes_6_out_ready; // @[pe.scala 268:49]
  assign PE_160_io_data_1_in_valid = PENetwork_25_io_to_pes_6_in_valid; // @[pe.scala 262:34]
  assign PE_160_io_data_1_in_bits = PENetwork_25_io_to_pes_6_in_bits; // @[pe.scala 262:34]
  assign PE_160_io_data_0_in_valid = PENetwork_6_io_to_pes_14_in_valid; // @[pe.scala 262:34]
  assign PE_160_io_data_0_in_bits = PENetwork_6_io_to_pes_14_in_bits; // @[pe.scala 262:34]
  assign PE_161_clock = clock;
  assign PE_161_reset = reset;
  assign PE_161_io_data_2_in_valid = PENetwork_40_io_to_pes_7_in_valid; // @[pe.scala 262:34]
  assign PE_161_io_data_2_in_bits = PENetwork_40_io_to_pes_7_in_bits; // @[pe.scala 262:34]
  assign PE_161_io_data_2_sig_stat2trans = PENetwork_40_io_to_pes_7_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_161_io_data_2_out_ready = PENetwork_40_io_to_pes_7_out_ready; // @[pe.scala 268:49]
  assign PE_161_io_data_1_in_valid = PENetwork_25_io_to_pes_7_in_valid; // @[pe.scala 262:34]
  assign PE_161_io_data_1_in_bits = PENetwork_25_io_to_pes_7_in_bits; // @[pe.scala 262:34]
  assign PE_161_io_data_0_in_valid = PENetwork_7_io_to_pes_14_in_valid; // @[pe.scala 262:34]
  assign PE_161_io_data_0_in_bits = PENetwork_7_io_to_pes_14_in_bits; // @[pe.scala 262:34]
  assign PE_162_clock = clock;
  assign PE_162_reset = reset;
  assign PE_162_io_data_2_in_valid = PENetwork_40_io_to_pes_8_in_valid; // @[pe.scala 262:34]
  assign PE_162_io_data_2_in_bits = PENetwork_40_io_to_pes_8_in_bits; // @[pe.scala 262:34]
  assign PE_162_io_data_2_sig_stat2trans = PENetwork_40_io_to_pes_8_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_162_io_data_2_out_ready = PENetwork_40_io_to_pes_8_out_ready; // @[pe.scala 268:49]
  assign PE_162_io_data_1_in_valid = PENetwork_25_io_to_pes_8_in_valid; // @[pe.scala 262:34]
  assign PE_162_io_data_1_in_bits = PENetwork_25_io_to_pes_8_in_bits; // @[pe.scala 262:34]
  assign PE_162_io_data_0_in_valid = PENetwork_8_io_to_pes_14_in_valid; // @[pe.scala 262:34]
  assign PE_162_io_data_0_in_bits = PENetwork_8_io_to_pes_14_in_bits; // @[pe.scala 262:34]
  assign PE_163_clock = clock;
  assign PE_163_reset = reset;
  assign PE_163_io_data_2_in_valid = PENetwork_40_io_to_pes_9_in_valid; // @[pe.scala 262:34]
  assign PE_163_io_data_2_in_bits = PENetwork_40_io_to_pes_9_in_bits; // @[pe.scala 262:34]
  assign PE_163_io_data_2_sig_stat2trans = PENetwork_40_io_to_pes_9_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_163_io_data_2_out_ready = PENetwork_40_io_to_pes_9_out_ready; // @[pe.scala 268:49]
  assign PE_163_io_data_1_in_valid = PENetwork_25_io_to_pes_9_in_valid; // @[pe.scala 262:34]
  assign PE_163_io_data_1_in_bits = PENetwork_25_io_to_pes_9_in_bits; // @[pe.scala 262:34]
  assign PE_163_io_data_0_in_valid = PENetwork_9_io_to_pes_14_in_valid; // @[pe.scala 262:34]
  assign PE_163_io_data_0_in_bits = PENetwork_9_io_to_pes_14_in_bits; // @[pe.scala 262:34]
  assign PE_164_clock = clock;
  assign PE_164_reset = reset;
  assign PE_164_io_data_2_in_valid = PENetwork_40_io_to_pes_10_in_valid; // @[pe.scala 262:34]
  assign PE_164_io_data_2_in_bits = PENetwork_40_io_to_pes_10_in_bits; // @[pe.scala 262:34]
  assign PE_164_io_data_2_sig_stat2trans = PENetwork_40_io_to_pes_10_sig_stat2trans; // @[pe.scala 265:52]
  assign PE_164_io_data_2_out_ready = 1'h1; // @[pe.scala 268:49]
  assign PE_164_io_data_1_in_valid = PENetwork_25_io_to_pes_10_in_valid; // @[pe.scala 262:34]
  assign PE_164_io_data_1_in_bits = PENetwork_25_io_to_pes_10_in_bits; // @[pe.scala 262:34]
  assign PE_164_io_data_0_in_valid = PENetwork_10_io_to_pes_14_in_valid; // @[pe.scala 262:34]
  assign PE_164_io_data_0_in_bits = PENetwork_10_io_to_pes_14_in_bits; // @[pe.scala 262:34]
  assign PENetwork_io_to_pes_0_out_valid = PE_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_io_to_pes_0_out_bits = PE_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_io_to_pes_1_out_valid = PE_11_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_io_to_pes_1_out_bits = PE_11_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_io_to_pes_2_out_valid = PE_22_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_io_to_pes_2_out_bits = PE_22_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_io_to_pes_3_out_valid = PE_33_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_io_to_pes_3_out_bits = PE_33_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_io_to_pes_4_out_valid = PE_44_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_io_to_pes_4_out_bits = PE_44_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_io_to_pes_5_out_valid = PE_55_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_io_to_pes_5_out_bits = PE_55_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_io_to_pes_6_out_valid = PE_66_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_io_to_pes_6_out_bits = PE_66_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_io_to_pes_7_out_valid = PE_77_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_io_to_pes_7_out_bits = PE_77_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_io_to_pes_8_out_valid = PE_88_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_io_to_pes_8_out_bits = PE_88_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_io_to_pes_9_out_valid = PE_99_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_io_to_pes_9_out_bits = PE_99_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_io_to_pes_10_out_valid = PE_110_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_io_to_pes_10_out_bits = PE_110_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_io_to_pes_11_out_valid = PE_121_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_io_to_pes_11_out_bits = PE_121_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_io_to_pes_12_out_valid = PE_132_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_io_to_pes_12_out_bits = PE_132_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_io_to_pes_13_out_valid = PE_143_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_io_to_pes_13_out_bits = PE_143_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_io_to_mem_valid = MemController_io_rd_data_valid; // @[pe.scala 315:29]
  assign PENetwork_io_to_mem_bits = MemController_io_rd_data_bits; // @[pe.scala 315:29]
  assign PENetwork_1_io_to_pes_0_out_valid = PE_1_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_1_io_to_pes_0_out_bits = PE_1_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_1_io_to_pes_1_out_valid = PE_12_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_1_io_to_pes_1_out_bits = PE_12_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_1_io_to_pes_2_out_valid = PE_23_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_1_io_to_pes_2_out_bits = PE_23_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_1_io_to_pes_3_out_valid = PE_34_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_1_io_to_pes_3_out_bits = PE_34_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_1_io_to_pes_4_out_valid = PE_45_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_1_io_to_pes_4_out_bits = PE_45_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_1_io_to_pes_5_out_valid = PE_56_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_1_io_to_pes_5_out_bits = PE_56_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_1_io_to_pes_6_out_valid = PE_67_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_1_io_to_pes_6_out_bits = PE_67_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_1_io_to_pes_7_out_valid = PE_78_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_1_io_to_pes_7_out_bits = PE_78_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_1_io_to_pes_8_out_valid = PE_89_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_1_io_to_pes_8_out_bits = PE_89_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_1_io_to_pes_9_out_valid = PE_100_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_1_io_to_pes_9_out_bits = PE_100_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_1_io_to_pes_10_out_valid = PE_111_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_1_io_to_pes_10_out_bits = PE_111_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_1_io_to_pes_11_out_valid = PE_122_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_1_io_to_pes_11_out_bits = PE_122_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_1_io_to_pes_12_out_valid = PE_133_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_1_io_to_pes_12_out_bits = PE_133_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_1_io_to_pes_13_out_valid = PE_144_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_1_io_to_pes_13_out_bits = PE_144_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_1_io_to_mem_valid = MemController_1_io_rd_data_valid; // @[pe.scala 315:29]
  assign PENetwork_1_io_to_mem_bits = MemController_1_io_rd_data_bits; // @[pe.scala 315:29]
  assign PENetwork_2_io_to_pes_0_out_valid = PE_2_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_2_io_to_pes_0_out_bits = PE_2_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_2_io_to_pes_1_out_valid = PE_13_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_2_io_to_pes_1_out_bits = PE_13_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_2_io_to_pes_2_out_valid = PE_24_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_2_io_to_pes_2_out_bits = PE_24_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_2_io_to_pes_3_out_valid = PE_35_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_2_io_to_pes_3_out_bits = PE_35_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_2_io_to_pes_4_out_valid = PE_46_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_2_io_to_pes_4_out_bits = PE_46_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_2_io_to_pes_5_out_valid = PE_57_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_2_io_to_pes_5_out_bits = PE_57_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_2_io_to_pes_6_out_valid = PE_68_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_2_io_to_pes_6_out_bits = PE_68_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_2_io_to_pes_7_out_valid = PE_79_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_2_io_to_pes_7_out_bits = PE_79_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_2_io_to_pes_8_out_valid = PE_90_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_2_io_to_pes_8_out_bits = PE_90_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_2_io_to_pes_9_out_valid = PE_101_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_2_io_to_pes_9_out_bits = PE_101_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_2_io_to_pes_10_out_valid = PE_112_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_2_io_to_pes_10_out_bits = PE_112_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_2_io_to_pes_11_out_valid = PE_123_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_2_io_to_pes_11_out_bits = PE_123_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_2_io_to_pes_12_out_valid = PE_134_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_2_io_to_pes_12_out_bits = PE_134_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_2_io_to_pes_13_out_valid = PE_145_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_2_io_to_pes_13_out_bits = PE_145_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_2_io_to_mem_valid = MemController_2_io_rd_data_valid; // @[pe.scala 315:29]
  assign PENetwork_2_io_to_mem_bits = MemController_2_io_rd_data_bits; // @[pe.scala 315:29]
  assign PENetwork_3_io_to_pes_0_out_valid = PE_3_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_3_io_to_pes_0_out_bits = PE_3_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_3_io_to_pes_1_out_valid = PE_14_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_3_io_to_pes_1_out_bits = PE_14_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_3_io_to_pes_2_out_valid = PE_25_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_3_io_to_pes_2_out_bits = PE_25_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_3_io_to_pes_3_out_valid = PE_36_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_3_io_to_pes_3_out_bits = PE_36_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_3_io_to_pes_4_out_valid = PE_47_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_3_io_to_pes_4_out_bits = PE_47_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_3_io_to_pes_5_out_valid = PE_58_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_3_io_to_pes_5_out_bits = PE_58_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_3_io_to_pes_6_out_valid = PE_69_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_3_io_to_pes_6_out_bits = PE_69_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_3_io_to_pes_7_out_valid = PE_80_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_3_io_to_pes_7_out_bits = PE_80_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_3_io_to_pes_8_out_valid = PE_91_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_3_io_to_pes_8_out_bits = PE_91_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_3_io_to_pes_9_out_valid = PE_102_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_3_io_to_pes_9_out_bits = PE_102_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_3_io_to_pes_10_out_valid = PE_113_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_3_io_to_pes_10_out_bits = PE_113_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_3_io_to_pes_11_out_valid = PE_124_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_3_io_to_pes_11_out_bits = PE_124_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_3_io_to_pes_12_out_valid = PE_135_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_3_io_to_pes_12_out_bits = PE_135_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_3_io_to_pes_13_out_valid = PE_146_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_3_io_to_pes_13_out_bits = PE_146_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_3_io_to_mem_valid = MemController_3_io_rd_data_valid; // @[pe.scala 315:29]
  assign PENetwork_3_io_to_mem_bits = MemController_3_io_rd_data_bits; // @[pe.scala 315:29]
  assign PENetwork_4_io_to_pes_0_out_valid = PE_4_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_4_io_to_pes_0_out_bits = PE_4_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_4_io_to_pes_1_out_valid = PE_15_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_4_io_to_pes_1_out_bits = PE_15_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_4_io_to_pes_2_out_valid = PE_26_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_4_io_to_pes_2_out_bits = PE_26_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_4_io_to_pes_3_out_valid = PE_37_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_4_io_to_pes_3_out_bits = PE_37_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_4_io_to_pes_4_out_valid = PE_48_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_4_io_to_pes_4_out_bits = PE_48_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_4_io_to_pes_5_out_valid = PE_59_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_4_io_to_pes_5_out_bits = PE_59_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_4_io_to_pes_6_out_valid = PE_70_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_4_io_to_pes_6_out_bits = PE_70_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_4_io_to_pes_7_out_valid = PE_81_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_4_io_to_pes_7_out_bits = PE_81_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_4_io_to_pes_8_out_valid = PE_92_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_4_io_to_pes_8_out_bits = PE_92_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_4_io_to_pes_9_out_valid = PE_103_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_4_io_to_pes_9_out_bits = PE_103_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_4_io_to_pes_10_out_valid = PE_114_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_4_io_to_pes_10_out_bits = PE_114_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_4_io_to_pes_11_out_valid = PE_125_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_4_io_to_pes_11_out_bits = PE_125_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_4_io_to_pes_12_out_valid = PE_136_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_4_io_to_pes_12_out_bits = PE_136_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_4_io_to_pes_13_out_valid = PE_147_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_4_io_to_pes_13_out_bits = PE_147_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_4_io_to_mem_valid = MemController_4_io_rd_data_valid; // @[pe.scala 315:29]
  assign PENetwork_4_io_to_mem_bits = MemController_4_io_rd_data_bits; // @[pe.scala 315:29]
  assign PENetwork_5_io_to_pes_0_out_valid = PE_5_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_5_io_to_pes_0_out_bits = PE_5_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_5_io_to_pes_1_out_valid = PE_16_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_5_io_to_pes_1_out_bits = PE_16_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_5_io_to_pes_2_out_valid = PE_27_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_5_io_to_pes_2_out_bits = PE_27_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_5_io_to_pes_3_out_valid = PE_38_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_5_io_to_pes_3_out_bits = PE_38_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_5_io_to_pes_4_out_valid = PE_49_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_5_io_to_pes_4_out_bits = PE_49_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_5_io_to_pes_5_out_valid = PE_60_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_5_io_to_pes_5_out_bits = PE_60_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_5_io_to_pes_6_out_valid = PE_71_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_5_io_to_pes_6_out_bits = PE_71_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_5_io_to_pes_7_out_valid = PE_82_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_5_io_to_pes_7_out_bits = PE_82_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_5_io_to_pes_8_out_valid = PE_93_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_5_io_to_pes_8_out_bits = PE_93_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_5_io_to_pes_9_out_valid = PE_104_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_5_io_to_pes_9_out_bits = PE_104_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_5_io_to_pes_10_out_valid = PE_115_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_5_io_to_pes_10_out_bits = PE_115_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_5_io_to_pes_11_out_valid = PE_126_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_5_io_to_pes_11_out_bits = PE_126_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_5_io_to_pes_12_out_valid = PE_137_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_5_io_to_pes_12_out_bits = PE_137_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_5_io_to_pes_13_out_valid = PE_148_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_5_io_to_pes_13_out_bits = PE_148_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_5_io_to_mem_valid = MemController_5_io_rd_data_valid; // @[pe.scala 315:29]
  assign PENetwork_5_io_to_mem_bits = MemController_5_io_rd_data_bits; // @[pe.scala 315:29]
  assign PENetwork_6_io_to_pes_0_out_valid = PE_6_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_6_io_to_pes_0_out_bits = PE_6_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_6_io_to_pes_1_out_valid = PE_17_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_6_io_to_pes_1_out_bits = PE_17_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_6_io_to_pes_2_out_valid = PE_28_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_6_io_to_pes_2_out_bits = PE_28_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_6_io_to_pes_3_out_valid = PE_39_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_6_io_to_pes_3_out_bits = PE_39_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_6_io_to_pes_4_out_valid = PE_50_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_6_io_to_pes_4_out_bits = PE_50_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_6_io_to_pes_5_out_valid = PE_61_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_6_io_to_pes_5_out_bits = PE_61_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_6_io_to_pes_6_out_valid = PE_72_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_6_io_to_pes_6_out_bits = PE_72_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_6_io_to_pes_7_out_valid = PE_83_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_6_io_to_pes_7_out_bits = PE_83_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_6_io_to_pes_8_out_valid = PE_94_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_6_io_to_pes_8_out_bits = PE_94_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_6_io_to_pes_9_out_valid = PE_105_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_6_io_to_pes_9_out_bits = PE_105_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_6_io_to_pes_10_out_valid = PE_116_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_6_io_to_pes_10_out_bits = PE_116_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_6_io_to_pes_11_out_valid = PE_127_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_6_io_to_pes_11_out_bits = PE_127_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_6_io_to_pes_12_out_valid = PE_138_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_6_io_to_pes_12_out_bits = PE_138_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_6_io_to_pes_13_out_valid = PE_149_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_6_io_to_pes_13_out_bits = PE_149_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_6_io_to_mem_valid = MemController_6_io_rd_data_valid; // @[pe.scala 315:29]
  assign PENetwork_6_io_to_mem_bits = MemController_6_io_rd_data_bits; // @[pe.scala 315:29]
  assign PENetwork_7_io_to_pes_0_out_valid = PE_7_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_7_io_to_pes_0_out_bits = PE_7_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_7_io_to_pes_1_out_valid = PE_18_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_7_io_to_pes_1_out_bits = PE_18_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_7_io_to_pes_2_out_valid = PE_29_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_7_io_to_pes_2_out_bits = PE_29_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_7_io_to_pes_3_out_valid = PE_40_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_7_io_to_pes_3_out_bits = PE_40_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_7_io_to_pes_4_out_valid = PE_51_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_7_io_to_pes_4_out_bits = PE_51_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_7_io_to_pes_5_out_valid = PE_62_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_7_io_to_pes_5_out_bits = PE_62_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_7_io_to_pes_6_out_valid = PE_73_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_7_io_to_pes_6_out_bits = PE_73_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_7_io_to_pes_7_out_valid = PE_84_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_7_io_to_pes_7_out_bits = PE_84_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_7_io_to_pes_8_out_valid = PE_95_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_7_io_to_pes_8_out_bits = PE_95_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_7_io_to_pes_9_out_valid = PE_106_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_7_io_to_pes_9_out_bits = PE_106_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_7_io_to_pes_10_out_valid = PE_117_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_7_io_to_pes_10_out_bits = PE_117_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_7_io_to_pes_11_out_valid = PE_128_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_7_io_to_pes_11_out_bits = PE_128_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_7_io_to_pes_12_out_valid = PE_139_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_7_io_to_pes_12_out_bits = PE_139_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_7_io_to_pes_13_out_valid = PE_150_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_7_io_to_pes_13_out_bits = PE_150_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_7_io_to_mem_valid = MemController_7_io_rd_data_valid; // @[pe.scala 315:29]
  assign PENetwork_7_io_to_mem_bits = MemController_7_io_rd_data_bits; // @[pe.scala 315:29]
  assign PENetwork_8_io_to_pes_0_out_valid = PE_8_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_8_io_to_pes_0_out_bits = PE_8_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_8_io_to_pes_1_out_valid = PE_19_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_8_io_to_pes_1_out_bits = PE_19_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_8_io_to_pes_2_out_valid = PE_30_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_8_io_to_pes_2_out_bits = PE_30_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_8_io_to_pes_3_out_valid = PE_41_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_8_io_to_pes_3_out_bits = PE_41_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_8_io_to_pes_4_out_valid = PE_52_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_8_io_to_pes_4_out_bits = PE_52_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_8_io_to_pes_5_out_valid = PE_63_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_8_io_to_pes_5_out_bits = PE_63_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_8_io_to_pes_6_out_valid = PE_74_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_8_io_to_pes_6_out_bits = PE_74_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_8_io_to_pes_7_out_valid = PE_85_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_8_io_to_pes_7_out_bits = PE_85_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_8_io_to_pes_8_out_valid = PE_96_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_8_io_to_pes_8_out_bits = PE_96_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_8_io_to_pes_9_out_valid = PE_107_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_8_io_to_pes_9_out_bits = PE_107_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_8_io_to_pes_10_out_valid = PE_118_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_8_io_to_pes_10_out_bits = PE_118_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_8_io_to_pes_11_out_valid = PE_129_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_8_io_to_pes_11_out_bits = PE_129_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_8_io_to_pes_12_out_valid = PE_140_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_8_io_to_pes_12_out_bits = PE_140_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_8_io_to_pes_13_out_valid = PE_151_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_8_io_to_pes_13_out_bits = PE_151_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_8_io_to_mem_valid = MemController_8_io_rd_data_valid; // @[pe.scala 315:29]
  assign PENetwork_8_io_to_mem_bits = MemController_8_io_rd_data_bits; // @[pe.scala 315:29]
  assign PENetwork_9_io_to_pes_0_out_valid = PE_9_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_9_io_to_pes_0_out_bits = PE_9_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_9_io_to_pes_1_out_valid = PE_20_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_9_io_to_pes_1_out_bits = PE_20_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_9_io_to_pes_2_out_valid = PE_31_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_9_io_to_pes_2_out_bits = PE_31_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_9_io_to_pes_3_out_valid = PE_42_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_9_io_to_pes_3_out_bits = PE_42_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_9_io_to_pes_4_out_valid = PE_53_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_9_io_to_pes_4_out_bits = PE_53_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_9_io_to_pes_5_out_valid = PE_64_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_9_io_to_pes_5_out_bits = PE_64_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_9_io_to_pes_6_out_valid = PE_75_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_9_io_to_pes_6_out_bits = PE_75_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_9_io_to_pes_7_out_valid = PE_86_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_9_io_to_pes_7_out_bits = PE_86_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_9_io_to_pes_8_out_valid = PE_97_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_9_io_to_pes_8_out_bits = PE_97_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_9_io_to_pes_9_out_valid = PE_108_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_9_io_to_pes_9_out_bits = PE_108_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_9_io_to_pes_10_out_valid = PE_119_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_9_io_to_pes_10_out_bits = PE_119_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_9_io_to_pes_11_out_valid = PE_130_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_9_io_to_pes_11_out_bits = PE_130_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_9_io_to_pes_12_out_valid = PE_141_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_9_io_to_pes_12_out_bits = PE_141_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_9_io_to_pes_13_out_valid = PE_152_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_9_io_to_pes_13_out_bits = PE_152_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_9_io_to_mem_valid = MemController_9_io_rd_data_valid; // @[pe.scala 315:29]
  assign PENetwork_9_io_to_mem_bits = MemController_9_io_rd_data_bits; // @[pe.scala 315:29]
  assign PENetwork_10_io_to_pes_0_out_valid = PE_10_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_10_io_to_pes_0_out_bits = PE_10_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_10_io_to_pes_1_out_valid = PE_21_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_10_io_to_pes_1_out_bits = PE_21_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_10_io_to_pes_2_out_valid = PE_32_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_10_io_to_pes_2_out_bits = PE_32_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_10_io_to_pes_3_out_valid = PE_43_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_10_io_to_pes_3_out_bits = PE_43_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_10_io_to_pes_4_out_valid = PE_54_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_10_io_to_pes_4_out_bits = PE_54_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_10_io_to_pes_5_out_valid = PE_65_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_10_io_to_pes_5_out_bits = PE_65_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_10_io_to_pes_6_out_valid = PE_76_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_10_io_to_pes_6_out_bits = PE_76_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_10_io_to_pes_7_out_valid = PE_87_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_10_io_to_pes_7_out_bits = PE_87_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_10_io_to_pes_8_out_valid = PE_98_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_10_io_to_pes_8_out_bits = PE_98_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_10_io_to_pes_9_out_valid = PE_109_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_10_io_to_pes_9_out_bits = PE_109_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_10_io_to_pes_10_out_valid = PE_120_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_10_io_to_pes_10_out_bits = PE_120_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_10_io_to_pes_11_out_valid = PE_131_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_10_io_to_pes_11_out_bits = PE_131_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_10_io_to_pes_12_out_valid = PE_142_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_10_io_to_pes_12_out_bits = PE_142_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_10_io_to_pes_13_out_valid = PE_153_io_data_0_out_valid; // @[pe.scala 261:36]
  assign PENetwork_10_io_to_pes_13_out_bits = PE_153_io_data_0_out_bits; // @[pe.scala 261:36]
  assign PENetwork_10_io_to_mem_valid = MemController_10_io_rd_data_valid; // @[pe.scala 315:29]
  assign PENetwork_10_io_to_mem_bits = MemController_10_io_rd_data_bits; // @[pe.scala 315:29]
  assign PENetwork_11_io_to_pes_0_out_valid = PE_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_11_io_to_pes_0_out_bits = PE_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_11_io_to_pes_1_out_valid = PE_1_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_11_io_to_pes_1_out_bits = PE_1_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_11_io_to_pes_2_out_valid = PE_2_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_11_io_to_pes_2_out_bits = PE_2_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_11_io_to_pes_3_out_valid = PE_3_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_11_io_to_pes_3_out_bits = PE_3_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_11_io_to_pes_4_out_valid = PE_4_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_11_io_to_pes_4_out_bits = PE_4_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_11_io_to_pes_5_out_valid = PE_5_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_11_io_to_pes_5_out_bits = PE_5_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_11_io_to_pes_6_out_valid = PE_6_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_11_io_to_pes_6_out_bits = PE_6_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_11_io_to_pes_7_out_valid = PE_7_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_11_io_to_pes_7_out_bits = PE_7_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_11_io_to_pes_8_out_valid = PE_8_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_11_io_to_pes_8_out_bits = PE_8_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_11_io_to_pes_9_out_valid = PE_9_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_11_io_to_pes_9_out_bits = PE_9_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_11_io_to_mem_valid = MemController_11_io_rd_data_valid; // @[pe.scala 315:29]
  assign PENetwork_11_io_to_mem_bits = MemController_11_io_rd_data_bits; // @[pe.scala 315:29]
  assign PENetwork_12_io_to_pes_0_out_valid = PE_11_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_12_io_to_pes_0_out_bits = PE_11_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_12_io_to_pes_1_out_valid = PE_12_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_12_io_to_pes_1_out_bits = PE_12_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_12_io_to_pes_2_out_valid = PE_13_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_12_io_to_pes_2_out_bits = PE_13_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_12_io_to_pes_3_out_valid = PE_14_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_12_io_to_pes_3_out_bits = PE_14_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_12_io_to_pes_4_out_valid = PE_15_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_12_io_to_pes_4_out_bits = PE_15_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_12_io_to_pes_5_out_valid = PE_16_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_12_io_to_pes_5_out_bits = PE_16_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_12_io_to_pes_6_out_valid = PE_17_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_12_io_to_pes_6_out_bits = PE_17_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_12_io_to_pes_7_out_valid = PE_18_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_12_io_to_pes_7_out_bits = PE_18_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_12_io_to_pes_8_out_valid = PE_19_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_12_io_to_pes_8_out_bits = PE_19_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_12_io_to_pes_9_out_valid = PE_20_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_12_io_to_pes_9_out_bits = PE_20_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_12_io_to_mem_valid = MemController_12_io_rd_data_valid; // @[pe.scala 315:29]
  assign PENetwork_12_io_to_mem_bits = MemController_12_io_rd_data_bits; // @[pe.scala 315:29]
  assign PENetwork_13_io_to_pes_0_out_valid = PE_22_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_13_io_to_pes_0_out_bits = PE_22_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_13_io_to_pes_1_out_valid = PE_23_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_13_io_to_pes_1_out_bits = PE_23_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_13_io_to_pes_2_out_valid = PE_24_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_13_io_to_pes_2_out_bits = PE_24_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_13_io_to_pes_3_out_valid = PE_25_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_13_io_to_pes_3_out_bits = PE_25_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_13_io_to_pes_4_out_valid = PE_26_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_13_io_to_pes_4_out_bits = PE_26_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_13_io_to_pes_5_out_valid = PE_27_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_13_io_to_pes_5_out_bits = PE_27_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_13_io_to_pes_6_out_valid = PE_28_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_13_io_to_pes_6_out_bits = PE_28_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_13_io_to_pes_7_out_valid = PE_29_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_13_io_to_pes_7_out_bits = PE_29_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_13_io_to_pes_8_out_valid = PE_30_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_13_io_to_pes_8_out_bits = PE_30_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_13_io_to_pes_9_out_valid = PE_31_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_13_io_to_pes_9_out_bits = PE_31_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_13_io_to_mem_valid = MemController_13_io_rd_data_valid; // @[pe.scala 315:29]
  assign PENetwork_13_io_to_mem_bits = MemController_13_io_rd_data_bits; // @[pe.scala 315:29]
  assign PENetwork_14_io_to_pes_0_out_valid = PE_33_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_14_io_to_pes_0_out_bits = PE_33_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_14_io_to_pes_1_out_valid = PE_34_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_14_io_to_pes_1_out_bits = PE_34_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_14_io_to_pes_2_out_valid = PE_35_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_14_io_to_pes_2_out_bits = PE_35_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_14_io_to_pes_3_out_valid = PE_36_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_14_io_to_pes_3_out_bits = PE_36_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_14_io_to_pes_4_out_valid = PE_37_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_14_io_to_pes_4_out_bits = PE_37_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_14_io_to_pes_5_out_valid = PE_38_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_14_io_to_pes_5_out_bits = PE_38_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_14_io_to_pes_6_out_valid = PE_39_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_14_io_to_pes_6_out_bits = PE_39_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_14_io_to_pes_7_out_valid = PE_40_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_14_io_to_pes_7_out_bits = PE_40_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_14_io_to_pes_8_out_valid = PE_41_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_14_io_to_pes_8_out_bits = PE_41_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_14_io_to_pes_9_out_valid = PE_42_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_14_io_to_pes_9_out_bits = PE_42_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_14_io_to_mem_valid = MemController_14_io_rd_data_valid; // @[pe.scala 315:29]
  assign PENetwork_14_io_to_mem_bits = MemController_14_io_rd_data_bits; // @[pe.scala 315:29]
  assign PENetwork_15_io_to_pes_0_out_valid = PE_44_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_15_io_to_pes_0_out_bits = PE_44_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_15_io_to_pes_1_out_valid = PE_45_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_15_io_to_pes_1_out_bits = PE_45_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_15_io_to_pes_2_out_valid = PE_46_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_15_io_to_pes_2_out_bits = PE_46_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_15_io_to_pes_3_out_valid = PE_47_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_15_io_to_pes_3_out_bits = PE_47_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_15_io_to_pes_4_out_valid = PE_48_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_15_io_to_pes_4_out_bits = PE_48_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_15_io_to_pes_5_out_valid = PE_49_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_15_io_to_pes_5_out_bits = PE_49_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_15_io_to_pes_6_out_valid = PE_50_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_15_io_to_pes_6_out_bits = PE_50_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_15_io_to_pes_7_out_valid = PE_51_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_15_io_to_pes_7_out_bits = PE_51_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_15_io_to_pes_8_out_valid = PE_52_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_15_io_to_pes_8_out_bits = PE_52_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_15_io_to_pes_9_out_valid = PE_53_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_15_io_to_pes_9_out_bits = PE_53_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_15_io_to_mem_valid = MemController_15_io_rd_data_valid; // @[pe.scala 315:29]
  assign PENetwork_15_io_to_mem_bits = MemController_15_io_rd_data_bits; // @[pe.scala 315:29]
  assign PENetwork_16_io_to_pes_0_out_valid = PE_55_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_16_io_to_pes_0_out_bits = PE_55_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_16_io_to_pes_1_out_valid = PE_56_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_16_io_to_pes_1_out_bits = PE_56_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_16_io_to_pes_2_out_valid = PE_57_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_16_io_to_pes_2_out_bits = PE_57_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_16_io_to_pes_3_out_valid = PE_58_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_16_io_to_pes_3_out_bits = PE_58_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_16_io_to_pes_4_out_valid = PE_59_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_16_io_to_pes_4_out_bits = PE_59_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_16_io_to_pes_5_out_valid = PE_60_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_16_io_to_pes_5_out_bits = PE_60_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_16_io_to_pes_6_out_valid = PE_61_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_16_io_to_pes_6_out_bits = PE_61_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_16_io_to_pes_7_out_valid = PE_62_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_16_io_to_pes_7_out_bits = PE_62_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_16_io_to_pes_8_out_valid = PE_63_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_16_io_to_pes_8_out_bits = PE_63_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_16_io_to_pes_9_out_valid = PE_64_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_16_io_to_pes_9_out_bits = PE_64_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_16_io_to_mem_valid = MemController_16_io_rd_data_valid; // @[pe.scala 315:29]
  assign PENetwork_16_io_to_mem_bits = MemController_16_io_rd_data_bits; // @[pe.scala 315:29]
  assign PENetwork_17_io_to_pes_0_out_valid = PE_66_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_17_io_to_pes_0_out_bits = PE_66_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_17_io_to_pes_1_out_valid = PE_67_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_17_io_to_pes_1_out_bits = PE_67_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_17_io_to_pes_2_out_valid = PE_68_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_17_io_to_pes_2_out_bits = PE_68_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_17_io_to_pes_3_out_valid = PE_69_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_17_io_to_pes_3_out_bits = PE_69_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_17_io_to_pes_4_out_valid = PE_70_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_17_io_to_pes_4_out_bits = PE_70_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_17_io_to_pes_5_out_valid = PE_71_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_17_io_to_pes_5_out_bits = PE_71_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_17_io_to_pes_6_out_valid = PE_72_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_17_io_to_pes_6_out_bits = PE_72_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_17_io_to_pes_7_out_valid = PE_73_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_17_io_to_pes_7_out_bits = PE_73_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_17_io_to_pes_8_out_valid = PE_74_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_17_io_to_pes_8_out_bits = PE_74_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_17_io_to_pes_9_out_valid = PE_75_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_17_io_to_pes_9_out_bits = PE_75_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_17_io_to_mem_valid = MemController_17_io_rd_data_valid; // @[pe.scala 315:29]
  assign PENetwork_17_io_to_mem_bits = MemController_17_io_rd_data_bits; // @[pe.scala 315:29]
  assign PENetwork_18_io_to_pes_0_out_valid = PE_77_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_18_io_to_pes_0_out_bits = PE_77_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_18_io_to_pes_1_out_valid = PE_78_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_18_io_to_pes_1_out_bits = PE_78_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_18_io_to_pes_2_out_valid = PE_79_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_18_io_to_pes_2_out_bits = PE_79_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_18_io_to_pes_3_out_valid = PE_80_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_18_io_to_pes_3_out_bits = PE_80_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_18_io_to_pes_4_out_valid = PE_81_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_18_io_to_pes_4_out_bits = PE_81_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_18_io_to_pes_5_out_valid = PE_82_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_18_io_to_pes_5_out_bits = PE_82_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_18_io_to_pes_6_out_valid = PE_83_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_18_io_to_pes_6_out_bits = PE_83_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_18_io_to_pes_7_out_valid = PE_84_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_18_io_to_pes_7_out_bits = PE_84_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_18_io_to_pes_8_out_valid = PE_85_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_18_io_to_pes_8_out_bits = PE_85_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_18_io_to_pes_9_out_valid = PE_86_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_18_io_to_pes_9_out_bits = PE_86_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_18_io_to_mem_valid = MemController_18_io_rd_data_valid; // @[pe.scala 315:29]
  assign PENetwork_18_io_to_mem_bits = MemController_18_io_rd_data_bits; // @[pe.scala 315:29]
  assign PENetwork_19_io_to_pes_0_out_valid = PE_88_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_19_io_to_pes_0_out_bits = PE_88_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_19_io_to_pes_1_out_valid = PE_89_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_19_io_to_pes_1_out_bits = PE_89_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_19_io_to_pes_2_out_valid = PE_90_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_19_io_to_pes_2_out_bits = PE_90_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_19_io_to_pes_3_out_valid = PE_91_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_19_io_to_pes_3_out_bits = PE_91_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_19_io_to_pes_4_out_valid = PE_92_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_19_io_to_pes_4_out_bits = PE_92_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_19_io_to_pes_5_out_valid = PE_93_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_19_io_to_pes_5_out_bits = PE_93_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_19_io_to_pes_6_out_valid = PE_94_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_19_io_to_pes_6_out_bits = PE_94_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_19_io_to_pes_7_out_valid = PE_95_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_19_io_to_pes_7_out_bits = PE_95_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_19_io_to_pes_8_out_valid = PE_96_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_19_io_to_pes_8_out_bits = PE_96_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_19_io_to_pes_9_out_valid = PE_97_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_19_io_to_pes_9_out_bits = PE_97_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_19_io_to_mem_valid = MemController_19_io_rd_data_valid; // @[pe.scala 315:29]
  assign PENetwork_19_io_to_mem_bits = MemController_19_io_rd_data_bits; // @[pe.scala 315:29]
  assign PENetwork_20_io_to_pes_0_out_valid = PE_99_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_20_io_to_pes_0_out_bits = PE_99_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_20_io_to_pes_1_out_valid = PE_100_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_20_io_to_pes_1_out_bits = PE_100_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_20_io_to_pes_2_out_valid = PE_101_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_20_io_to_pes_2_out_bits = PE_101_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_20_io_to_pes_3_out_valid = PE_102_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_20_io_to_pes_3_out_bits = PE_102_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_20_io_to_pes_4_out_valid = PE_103_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_20_io_to_pes_4_out_bits = PE_103_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_20_io_to_pes_5_out_valid = PE_104_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_20_io_to_pes_5_out_bits = PE_104_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_20_io_to_pes_6_out_valid = PE_105_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_20_io_to_pes_6_out_bits = PE_105_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_20_io_to_pes_7_out_valid = PE_106_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_20_io_to_pes_7_out_bits = PE_106_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_20_io_to_pes_8_out_valid = PE_107_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_20_io_to_pes_8_out_bits = PE_107_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_20_io_to_pes_9_out_valid = PE_108_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_20_io_to_pes_9_out_bits = PE_108_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_20_io_to_mem_valid = MemController_20_io_rd_data_valid; // @[pe.scala 315:29]
  assign PENetwork_20_io_to_mem_bits = MemController_20_io_rd_data_bits; // @[pe.scala 315:29]
  assign PENetwork_21_io_to_pes_0_out_valid = PE_110_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_21_io_to_pes_0_out_bits = PE_110_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_21_io_to_pes_1_out_valid = PE_111_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_21_io_to_pes_1_out_bits = PE_111_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_21_io_to_pes_2_out_valid = PE_112_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_21_io_to_pes_2_out_bits = PE_112_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_21_io_to_pes_3_out_valid = PE_113_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_21_io_to_pes_3_out_bits = PE_113_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_21_io_to_pes_4_out_valid = PE_114_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_21_io_to_pes_4_out_bits = PE_114_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_21_io_to_pes_5_out_valid = PE_115_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_21_io_to_pes_5_out_bits = PE_115_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_21_io_to_pes_6_out_valid = PE_116_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_21_io_to_pes_6_out_bits = PE_116_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_21_io_to_pes_7_out_valid = PE_117_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_21_io_to_pes_7_out_bits = PE_117_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_21_io_to_pes_8_out_valid = PE_118_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_21_io_to_pes_8_out_bits = PE_118_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_21_io_to_pes_9_out_valid = PE_119_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_21_io_to_pes_9_out_bits = PE_119_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_21_io_to_mem_valid = MemController_21_io_rd_data_valid; // @[pe.scala 315:29]
  assign PENetwork_21_io_to_mem_bits = MemController_21_io_rd_data_bits; // @[pe.scala 315:29]
  assign PENetwork_22_io_to_pes_0_out_valid = PE_121_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_22_io_to_pes_0_out_bits = PE_121_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_22_io_to_pes_1_out_valid = PE_122_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_22_io_to_pes_1_out_bits = PE_122_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_22_io_to_pes_2_out_valid = PE_123_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_22_io_to_pes_2_out_bits = PE_123_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_22_io_to_pes_3_out_valid = PE_124_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_22_io_to_pes_3_out_bits = PE_124_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_22_io_to_pes_4_out_valid = PE_125_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_22_io_to_pes_4_out_bits = PE_125_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_22_io_to_pes_5_out_valid = PE_126_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_22_io_to_pes_5_out_bits = PE_126_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_22_io_to_pes_6_out_valid = PE_127_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_22_io_to_pes_6_out_bits = PE_127_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_22_io_to_pes_7_out_valid = PE_128_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_22_io_to_pes_7_out_bits = PE_128_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_22_io_to_pes_8_out_valid = PE_129_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_22_io_to_pes_8_out_bits = PE_129_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_22_io_to_pes_9_out_valid = PE_130_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_22_io_to_pes_9_out_bits = PE_130_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_22_io_to_mem_valid = MemController_22_io_rd_data_valid; // @[pe.scala 315:29]
  assign PENetwork_22_io_to_mem_bits = MemController_22_io_rd_data_bits; // @[pe.scala 315:29]
  assign PENetwork_23_io_to_pes_0_out_valid = PE_132_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_23_io_to_pes_0_out_bits = PE_132_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_23_io_to_pes_1_out_valid = PE_133_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_23_io_to_pes_1_out_bits = PE_133_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_23_io_to_pes_2_out_valid = PE_134_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_23_io_to_pes_2_out_bits = PE_134_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_23_io_to_pes_3_out_valid = PE_135_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_23_io_to_pes_3_out_bits = PE_135_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_23_io_to_pes_4_out_valid = PE_136_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_23_io_to_pes_4_out_bits = PE_136_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_23_io_to_pes_5_out_valid = PE_137_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_23_io_to_pes_5_out_bits = PE_137_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_23_io_to_pes_6_out_valid = PE_138_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_23_io_to_pes_6_out_bits = PE_138_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_23_io_to_pes_7_out_valid = PE_139_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_23_io_to_pes_7_out_bits = PE_139_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_23_io_to_pes_8_out_valid = PE_140_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_23_io_to_pes_8_out_bits = PE_140_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_23_io_to_pes_9_out_valid = PE_141_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_23_io_to_pes_9_out_bits = PE_141_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_23_io_to_mem_valid = MemController_23_io_rd_data_valid; // @[pe.scala 315:29]
  assign PENetwork_23_io_to_mem_bits = MemController_23_io_rd_data_bits; // @[pe.scala 315:29]
  assign PENetwork_24_io_to_pes_0_out_valid = PE_143_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_24_io_to_pes_0_out_bits = PE_143_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_24_io_to_pes_1_out_valid = PE_144_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_24_io_to_pes_1_out_bits = PE_144_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_24_io_to_pes_2_out_valid = PE_145_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_24_io_to_pes_2_out_bits = PE_145_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_24_io_to_pes_3_out_valid = PE_146_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_24_io_to_pes_3_out_bits = PE_146_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_24_io_to_pes_4_out_valid = PE_147_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_24_io_to_pes_4_out_bits = PE_147_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_24_io_to_pes_5_out_valid = PE_148_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_24_io_to_pes_5_out_bits = PE_148_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_24_io_to_pes_6_out_valid = PE_149_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_24_io_to_pes_6_out_bits = PE_149_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_24_io_to_pes_7_out_valid = PE_150_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_24_io_to_pes_7_out_bits = PE_150_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_24_io_to_pes_8_out_valid = PE_151_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_24_io_to_pes_8_out_bits = PE_151_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_24_io_to_pes_9_out_valid = PE_152_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_24_io_to_pes_9_out_bits = PE_152_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_24_io_to_mem_valid = MemController_24_io_rd_data_valid; // @[pe.scala 315:29]
  assign PENetwork_24_io_to_mem_bits = MemController_24_io_rd_data_bits; // @[pe.scala 315:29]
  assign PENetwork_25_io_to_pes_0_out_valid = PE_154_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_25_io_to_pes_0_out_bits = PE_154_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_25_io_to_pes_1_out_valid = PE_155_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_25_io_to_pes_1_out_bits = PE_155_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_25_io_to_pes_2_out_valid = PE_156_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_25_io_to_pes_2_out_bits = PE_156_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_25_io_to_pes_3_out_valid = PE_157_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_25_io_to_pes_3_out_bits = PE_157_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_25_io_to_pes_4_out_valid = PE_158_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_25_io_to_pes_4_out_bits = PE_158_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_25_io_to_pes_5_out_valid = PE_159_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_25_io_to_pes_5_out_bits = PE_159_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_25_io_to_pes_6_out_valid = PE_160_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_25_io_to_pes_6_out_bits = PE_160_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_25_io_to_pes_7_out_valid = PE_161_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_25_io_to_pes_7_out_bits = PE_161_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_25_io_to_pes_8_out_valid = PE_162_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_25_io_to_pes_8_out_bits = PE_162_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_25_io_to_pes_9_out_valid = PE_163_io_data_1_out_valid; // @[pe.scala 261:36]
  assign PENetwork_25_io_to_pes_9_out_bits = PE_163_io_data_1_out_bits; // @[pe.scala 261:36]
  assign PENetwork_25_io_to_mem_valid = MemController_25_io_rd_data_valid; // @[pe.scala 315:29]
  assign PENetwork_25_io_to_mem_bits = MemController_25_io_rd_data_bits; // @[pe.scala 315:29]
  assign PENetwork_26_clock = clock;
  assign PENetwork_26_io_to_pes_0_out_valid = PE_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_26_io_to_pes_0_out_bits = PE_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_26_io_to_pes_1_out_valid = PE_1_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_26_io_to_pes_1_out_bits = PE_1_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_26_io_to_pes_1_in_ready = PE_1_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_26_io_to_pes_2_out_valid = PE_2_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_26_io_to_pes_2_out_bits = PE_2_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_26_io_to_pes_2_in_ready = PE_2_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_26_io_to_pes_3_out_valid = PE_3_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_26_io_to_pes_3_out_bits = PE_3_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_26_io_to_pes_3_in_ready = PE_3_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_26_io_to_pes_4_out_valid = PE_4_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_26_io_to_pes_4_out_bits = PE_4_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_26_io_to_pes_4_in_ready = PE_4_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_26_io_to_pes_5_out_valid = PE_5_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_26_io_to_pes_5_out_bits = PE_5_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_26_io_to_pes_5_in_ready = PE_5_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_26_io_to_pes_6_out_valid = PE_6_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_26_io_to_pes_6_out_bits = PE_6_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_26_io_to_pes_6_in_ready = PE_6_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_26_io_to_pes_7_out_valid = PE_7_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_26_io_to_pes_7_out_bits = PE_7_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_26_io_to_pes_7_in_ready = PE_7_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_26_io_to_pes_8_out_valid = PE_8_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_26_io_to_pes_8_out_bits = PE_8_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_26_io_to_pes_8_in_ready = PE_8_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_26_io_to_pes_9_out_valid = PE_9_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_26_io_to_pes_9_out_bits = PE_9_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_26_io_to_pes_9_in_ready = PE_9_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_26_io_to_pes_10_out_valid = PE_10_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_26_io_to_pes_10_out_bits = PE_10_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_26_io_to_pes_10_in_ready = PE_10_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_26_io_sig_stat2trans = MultiDimTime_io_index_1 == 16'h0; // @[pe.scala 281:43]
  assign PENetwork_27_clock = clock;
  assign PENetwork_27_io_to_pes_0_out_valid = PE_11_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_27_io_to_pes_0_out_bits = PE_11_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_27_io_to_pes_1_out_valid = PE_12_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_27_io_to_pes_1_out_bits = PE_12_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_27_io_to_pes_1_in_ready = PE_12_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_27_io_to_pes_2_out_valid = PE_13_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_27_io_to_pes_2_out_bits = PE_13_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_27_io_to_pes_2_in_ready = PE_13_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_27_io_to_pes_3_out_valid = PE_14_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_27_io_to_pes_3_out_bits = PE_14_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_27_io_to_pes_3_in_ready = PE_14_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_27_io_to_pes_4_out_valid = PE_15_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_27_io_to_pes_4_out_bits = PE_15_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_27_io_to_pes_4_in_ready = PE_15_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_27_io_to_pes_5_out_valid = PE_16_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_27_io_to_pes_5_out_bits = PE_16_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_27_io_to_pes_5_in_ready = PE_16_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_27_io_to_pes_6_out_valid = PE_17_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_27_io_to_pes_6_out_bits = PE_17_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_27_io_to_pes_6_in_ready = PE_17_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_27_io_to_pes_7_out_valid = PE_18_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_27_io_to_pes_7_out_bits = PE_18_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_27_io_to_pes_7_in_ready = PE_18_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_27_io_to_pes_8_out_valid = PE_19_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_27_io_to_pes_8_out_bits = PE_19_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_27_io_to_pes_8_in_ready = PE_19_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_27_io_to_pes_9_out_valid = PE_20_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_27_io_to_pes_9_out_bits = PE_20_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_27_io_to_pes_9_in_ready = PE_20_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_27_io_to_pes_10_out_valid = PE_21_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_27_io_to_pes_10_out_bits = PE_21_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_27_io_to_pes_10_in_ready = PE_21_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_27_io_sig_stat2trans = MultiDimTime_io_index_1 == 16'h0; // @[pe.scala 281:43]
  assign PENetwork_28_clock = clock;
  assign PENetwork_28_io_to_pes_0_out_valid = PE_22_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_28_io_to_pes_0_out_bits = PE_22_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_28_io_to_pes_1_out_valid = PE_23_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_28_io_to_pes_1_out_bits = PE_23_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_28_io_to_pes_1_in_ready = PE_23_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_28_io_to_pes_2_out_valid = PE_24_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_28_io_to_pes_2_out_bits = PE_24_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_28_io_to_pes_2_in_ready = PE_24_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_28_io_to_pes_3_out_valid = PE_25_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_28_io_to_pes_3_out_bits = PE_25_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_28_io_to_pes_3_in_ready = PE_25_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_28_io_to_pes_4_out_valid = PE_26_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_28_io_to_pes_4_out_bits = PE_26_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_28_io_to_pes_4_in_ready = PE_26_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_28_io_to_pes_5_out_valid = PE_27_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_28_io_to_pes_5_out_bits = PE_27_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_28_io_to_pes_5_in_ready = PE_27_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_28_io_to_pes_6_out_valid = PE_28_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_28_io_to_pes_6_out_bits = PE_28_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_28_io_to_pes_6_in_ready = PE_28_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_28_io_to_pes_7_out_valid = PE_29_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_28_io_to_pes_7_out_bits = PE_29_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_28_io_to_pes_7_in_ready = PE_29_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_28_io_to_pes_8_out_valid = PE_30_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_28_io_to_pes_8_out_bits = PE_30_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_28_io_to_pes_8_in_ready = PE_30_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_28_io_to_pes_9_out_valid = PE_31_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_28_io_to_pes_9_out_bits = PE_31_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_28_io_to_pes_9_in_ready = PE_31_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_28_io_to_pes_10_out_valid = PE_32_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_28_io_to_pes_10_out_bits = PE_32_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_28_io_to_pes_10_in_ready = PE_32_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_28_io_sig_stat2trans = MultiDimTime_io_index_1 == 16'h0; // @[pe.scala 281:43]
  assign PENetwork_29_clock = clock;
  assign PENetwork_29_io_to_pes_0_out_valid = PE_33_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_29_io_to_pes_0_out_bits = PE_33_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_29_io_to_pes_1_out_valid = PE_34_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_29_io_to_pes_1_out_bits = PE_34_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_29_io_to_pes_1_in_ready = PE_34_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_29_io_to_pes_2_out_valid = PE_35_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_29_io_to_pes_2_out_bits = PE_35_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_29_io_to_pes_2_in_ready = PE_35_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_29_io_to_pes_3_out_valid = PE_36_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_29_io_to_pes_3_out_bits = PE_36_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_29_io_to_pes_3_in_ready = PE_36_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_29_io_to_pes_4_out_valid = PE_37_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_29_io_to_pes_4_out_bits = PE_37_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_29_io_to_pes_4_in_ready = PE_37_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_29_io_to_pes_5_out_valid = PE_38_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_29_io_to_pes_5_out_bits = PE_38_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_29_io_to_pes_5_in_ready = PE_38_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_29_io_to_pes_6_out_valid = PE_39_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_29_io_to_pes_6_out_bits = PE_39_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_29_io_to_pes_6_in_ready = PE_39_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_29_io_to_pes_7_out_valid = PE_40_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_29_io_to_pes_7_out_bits = PE_40_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_29_io_to_pes_7_in_ready = PE_40_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_29_io_to_pes_8_out_valid = PE_41_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_29_io_to_pes_8_out_bits = PE_41_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_29_io_to_pes_8_in_ready = PE_41_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_29_io_to_pes_9_out_valid = PE_42_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_29_io_to_pes_9_out_bits = PE_42_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_29_io_to_pes_9_in_ready = PE_42_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_29_io_to_pes_10_out_valid = PE_43_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_29_io_to_pes_10_out_bits = PE_43_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_29_io_to_pes_10_in_ready = PE_43_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_29_io_sig_stat2trans = MultiDimTime_io_index_1 == 16'h0; // @[pe.scala 281:43]
  assign PENetwork_30_clock = clock;
  assign PENetwork_30_io_to_pes_0_out_valid = PE_44_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_30_io_to_pes_0_out_bits = PE_44_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_30_io_to_pes_1_out_valid = PE_45_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_30_io_to_pes_1_out_bits = PE_45_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_30_io_to_pes_1_in_ready = PE_45_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_30_io_to_pes_2_out_valid = PE_46_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_30_io_to_pes_2_out_bits = PE_46_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_30_io_to_pes_2_in_ready = PE_46_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_30_io_to_pes_3_out_valid = PE_47_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_30_io_to_pes_3_out_bits = PE_47_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_30_io_to_pes_3_in_ready = PE_47_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_30_io_to_pes_4_out_valid = PE_48_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_30_io_to_pes_4_out_bits = PE_48_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_30_io_to_pes_4_in_ready = PE_48_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_30_io_to_pes_5_out_valid = PE_49_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_30_io_to_pes_5_out_bits = PE_49_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_30_io_to_pes_5_in_ready = PE_49_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_30_io_to_pes_6_out_valid = PE_50_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_30_io_to_pes_6_out_bits = PE_50_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_30_io_to_pes_6_in_ready = PE_50_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_30_io_to_pes_7_out_valid = PE_51_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_30_io_to_pes_7_out_bits = PE_51_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_30_io_to_pes_7_in_ready = PE_51_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_30_io_to_pes_8_out_valid = PE_52_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_30_io_to_pes_8_out_bits = PE_52_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_30_io_to_pes_8_in_ready = PE_52_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_30_io_to_pes_9_out_valid = PE_53_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_30_io_to_pes_9_out_bits = PE_53_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_30_io_to_pes_9_in_ready = PE_53_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_30_io_to_pes_10_out_valid = PE_54_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_30_io_to_pes_10_out_bits = PE_54_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_30_io_to_pes_10_in_ready = PE_54_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_30_io_sig_stat2trans = MultiDimTime_io_index_1 == 16'h0; // @[pe.scala 281:43]
  assign PENetwork_31_clock = clock;
  assign PENetwork_31_io_to_pes_0_out_valid = PE_55_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_31_io_to_pes_0_out_bits = PE_55_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_31_io_to_pes_1_out_valid = PE_56_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_31_io_to_pes_1_out_bits = PE_56_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_31_io_to_pes_1_in_ready = PE_56_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_31_io_to_pes_2_out_valid = PE_57_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_31_io_to_pes_2_out_bits = PE_57_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_31_io_to_pes_2_in_ready = PE_57_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_31_io_to_pes_3_out_valid = PE_58_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_31_io_to_pes_3_out_bits = PE_58_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_31_io_to_pes_3_in_ready = PE_58_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_31_io_to_pes_4_out_valid = PE_59_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_31_io_to_pes_4_out_bits = PE_59_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_31_io_to_pes_4_in_ready = PE_59_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_31_io_to_pes_5_out_valid = PE_60_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_31_io_to_pes_5_out_bits = PE_60_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_31_io_to_pes_5_in_ready = PE_60_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_31_io_to_pes_6_out_valid = PE_61_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_31_io_to_pes_6_out_bits = PE_61_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_31_io_to_pes_6_in_ready = PE_61_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_31_io_to_pes_7_out_valid = PE_62_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_31_io_to_pes_7_out_bits = PE_62_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_31_io_to_pes_7_in_ready = PE_62_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_31_io_to_pes_8_out_valid = PE_63_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_31_io_to_pes_8_out_bits = PE_63_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_31_io_to_pes_8_in_ready = PE_63_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_31_io_to_pes_9_out_valid = PE_64_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_31_io_to_pes_9_out_bits = PE_64_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_31_io_to_pes_9_in_ready = PE_64_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_31_io_to_pes_10_out_valid = PE_65_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_31_io_to_pes_10_out_bits = PE_65_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_31_io_to_pes_10_in_ready = PE_65_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_31_io_sig_stat2trans = MultiDimTime_io_index_1 == 16'h0; // @[pe.scala 281:43]
  assign PENetwork_32_clock = clock;
  assign PENetwork_32_io_to_pes_0_out_valid = PE_66_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_32_io_to_pes_0_out_bits = PE_66_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_32_io_to_pes_1_out_valid = PE_67_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_32_io_to_pes_1_out_bits = PE_67_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_32_io_to_pes_1_in_ready = PE_67_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_32_io_to_pes_2_out_valid = PE_68_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_32_io_to_pes_2_out_bits = PE_68_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_32_io_to_pes_2_in_ready = PE_68_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_32_io_to_pes_3_out_valid = PE_69_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_32_io_to_pes_3_out_bits = PE_69_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_32_io_to_pes_3_in_ready = PE_69_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_32_io_to_pes_4_out_valid = PE_70_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_32_io_to_pes_4_out_bits = PE_70_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_32_io_to_pes_4_in_ready = PE_70_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_32_io_to_pes_5_out_valid = PE_71_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_32_io_to_pes_5_out_bits = PE_71_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_32_io_to_pes_5_in_ready = PE_71_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_32_io_to_pes_6_out_valid = PE_72_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_32_io_to_pes_6_out_bits = PE_72_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_32_io_to_pes_6_in_ready = PE_72_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_32_io_to_pes_7_out_valid = PE_73_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_32_io_to_pes_7_out_bits = PE_73_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_32_io_to_pes_7_in_ready = PE_73_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_32_io_to_pes_8_out_valid = PE_74_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_32_io_to_pes_8_out_bits = PE_74_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_32_io_to_pes_8_in_ready = PE_74_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_32_io_to_pes_9_out_valid = PE_75_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_32_io_to_pes_9_out_bits = PE_75_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_32_io_to_pes_9_in_ready = PE_75_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_32_io_to_pes_10_out_valid = PE_76_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_32_io_to_pes_10_out_bits = PE_76_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_32_io_to_pes_10_in_ready = PE_76_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_32_io_sig_stat2trans = MultiDimTime_io_index_1 == 16'h0; // @[pe.scala 281:43]
  assign PENetwork_33_clock = clock;
  assign PENetwork_33_io_to_pes_0_out_valid = PE_77_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_33_io_to_pes_0_out_bits = PE_77_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_33_io_to_pes_1_out_valid = PE_78_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_33_io_to_pes_1_out_bits = PE_78_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_33_io_to_pes_1_in_ready = PE_78_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_33_io_to_pes_2_out_valid = PE_79_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_33_io_to_pes_2_out_bits = PE_79_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_33_io_to_pes_2_in_ready = PE_79_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_33_io_to_pes_3_out_valid = PE_80_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_33_io_to_pes_3_out_bits = PE_80_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_33_io_to_pes_3_in_ready = PE_80_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_33_io_to_pes_4_out_valid = PE_81_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_33_io_to_pes_4_out_bits = PE_81_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_33_io_to_pes_4_in_ready = PE_81_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_33_io_to_pes_5_out_valid = PE_82_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_33_io_to_pes_5_out_bits = PE_82_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_33_io_to_pes_5_in_ready = PE_82_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_33_io_to_pes_6_out_valid = PE_83_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_33_io_to_pes_6_out_bits = PE_83_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_33_io_to_pes_6_in_ready = PE_83_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_33_io_to_pes_7_out_valid = PE_84_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_33_io_to_pes_7_out_bits = PE_84_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_33_io_to_pes_7_in_ready = PE_84_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_33_io_to_pes_8_out_valid = PE_85_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_33_io_to_pes_8_out_bits = PE_85_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_33_io_to_pes_8_in_ready = PE_85_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_33_io_to_pes_9_out_valid = PE_86_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_33_io_to_pes_9_out_bits = PE_86_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_33_io_to_pes_9_in_ready = PE_86_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_33_io_to_pes_10_out_valid = PE_87_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_33_io_to_pes_10_out_bits = PE_87_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_33_io_to_pes_10_in_ready = PE_87_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_33_io_sig_stat2trans = MultiDimTime_io_index_1 == 16'h0; // @[pe.scala 281:43]
  assign PENetwork_34_clock = clock;
  assign PENetwork_34_io_to_pes_0_out_valid = PE_88_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_34_io_to_pes_0_out_bits = PE_88_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_34_io_to_pes_1_out_valid = PE_89_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_34_io_to_pes_1_out_bits = PE_89_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_34_io_to_pes_1_in_ready = PE_89_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_34_io_to_pes_2_out_valid = PE_90_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_34_io_to_pes_2_out_bits = PE_90_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_34_io_to_pes_2_in_ready = PE_90_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_34_io_to_pes_3_out_valid = PE_91_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_34_io_to_pes_3_out_bits = PE_91_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_34_io_to_pes_3_in_ready = PE_91_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_34_io_to_pes_4_out_valid = PE_92_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_34_io_to_pes_4_out_bits = PE_92_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_34_io_to_pes_4_in_ready = PE_92_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_34_io_to_pes_5_out_valid = PE_93_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_34_io_to_pes_5_out_bits = PE_93_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_34_io_to_pes_5_in_ready = PE_93_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_34_io_to_pes_6_out_valid = PE_94_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_34_io_to_pes_6_out_bits = PE_94_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_34_io_to_pes_6_in_ready = PE_94_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_34_io_to_pes_7_out_valid = PE_95_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_34_io_to_pes_7_out_bits = PE_95_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_34_io_to_pes_7_in_ready = PE_95_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_34_io_to_pes_8_out_valid = PE_96_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_34_io_to_pes_8_out_bits = PE_96_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_34_io_to_pes_8_in_ready = PE_96_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_34_io_to_pes_9_out_valid = PE_97_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_34_io_to_pes_9_out_bits = PE_97_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_34_io_to_pes_9_in_ready = PE_97_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_34_io_to_pes_10_out_valid = PE_98_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_34_io_to_pes_10_out_bits = PE_98_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_34_io_to_pes_10_in_ready = PE_98_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_34_io_sig_stat2trans = MultiDimTime_io_index_1 == 16'h0; // @[pe.scala 281:43]
  assign PENetwork_35_clock = clock;
  assign PENetwork_35_io_to_pes_0_out_valid = PE_99_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_35_io_to_pes_0_out_bits = PE_99_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_35_io_to_pes_1_out_valid = PE_100_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_35_io_to_pes_1_out_bits = PE_100_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_35_io_to_pes_1_in_ready = PE_100_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_35_io_to_pes_2_out_valid = PE_101_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_35_io_to_pes_2_out_bits = PE_101_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_35_io_to_pes_2_in_ready = PE_101_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_35_io_to_pes_3_out_valid = PE_102_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_35_io_to_pes_3_out_bits = PE_102_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_35_io_to_pes_3_in_ready = PE_102_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_35_io_to_pes_4_out_valid = PE_103_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_35_io_to_pes_4_out_bits = PE_103_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_35_io_to_pes_4_in_ready = PE_103_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_35_io_to_pes_5_out_valid = PE_104_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_35_io_to_pes_5_out_bits = PE_104_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_35_io_to_pes_5_in_ready = PE_104_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_35_io_to_pes_6_out_valid = PE_105_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_35_io_to_pes_6_out_bits = PE_105_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_35_io_to_pes_6_in_ready = PE_105_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_35_io_to_pes_7_out_valid = PE_106_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_35_io_to_pes_7_out_bits = PE_106_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_35_io_to_pes_7_in_ready = PE_106_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_35_io_to_pes_8_out_valid = PE_107_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_35_io_to_pes_8_out_bits = PE_107_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_35_io_to_pes_8_in_ready = PE_107_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_35_io_to_pes_9_out_valid = PE_108_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_35_io_to_pes_9_out_bits = PE_108_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_35_io_to_pes_9_in_ready = PE_108_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_35_io_to_pes_10_out_valid = PE_109_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_35_io_to_pes_10_out_bits = PE_109_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_35_io_to_pes_10_in_ready = PE_109_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_35_io_sig_stat2trans = MultiDimTime_io_index_1 == 16'h0; // @[pe.scala 281:43]
  assign PENetwork_36_clock = clock;
  assign PENetwork_36_io_to_pes_0_out_valid = PE_110_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_36_io_to_pes_0_out_bits = PE_110_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_36_io_to_pes_1_out_valid = PE_111_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_36_io_to_pes_1_out_bits = PE_111_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_36_io_to_pes_1_in_ready = PE_111_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_36_io_to_pes_2_out_valid = PE_112_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_36_io_to_pes_2_out_bits = PE_112_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_36_io_to_pes_2_in_ready = PE_112_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_36_io_to_pes_3_out_valid = PE_113_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_36_io_to_pes_3_out_bits = PE_113_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_36_io_to_pes_3_in_ready = PE_113_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_36_io_to_pes_4_out_valid = PE_114_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_36_io_to_pes_4_out_bits = PE_114_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_36_io_to_pes_4_in_ready = PE_114_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_36_io_to_pes_5_out_valid = PE_115_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_36_io_to_pes_5_out_bits = PE_115_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_36_io_to_pes_5_in_ready = PE_115_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_36_io_to_pes_6_out_valid = PE_116_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_36_io_to_pes_6_out_bits = PE_116_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_36_io_to_pes_6_in_ready = PE_116_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_36_io_to_pes_7_out_valid = PE_117_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_36_io_to_pes_7_out_bits = PE_117_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_36_io_to_pes_7_in_ready = PE_117_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_36_io_to_pes_8_out_valid = PE_118_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_36_io_to_pes_8_out_bits = PE_118_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_36_io_to_pes_8_in_ready = PE_118_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_36_io_to_pes_9_out_valid = PE_119_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_36_io_to_pes_9_out_bits = PE_119_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_36_io_to_pes_9_in_ready = PE_119_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_36_io_to_pes_10_out_valid = PE_120_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_36_io_to_pes_10_out_bits = PE_120_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_36_io_to_pes_10_in_ready = PE_120_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_36_io_sig_stat2trans = MultiDimTime_io_index_1 == 16'h0; // @[pe.scala 281:43]
  assign PENetwork_37_clock = clock;
  assign PENetwork_37_io_to_pes_0_out_valid = PE_121_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_37_io_to_pes_0_out_bits = PE_121_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_37_io_to_pes_1_out_valid = PE_122_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_37_io_to_pes_1_out_bits = PE_122_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_37_io_to_pes_1_in_ready = PE_122_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_37_io_to_pes_2_out_valid = PE_123_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_37_io_to_pes_2_out_bits = PE_123_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_37_io_to_pes_2_in_ready = PE_123_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_37_io_to_pes_3_out_valid = PE_124_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_37_io_to_pes_3_out_bits = PE_124_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_37_io_to_pes_3_in_ready = PE_124_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_37_io_to_pes_4_out_valid = PE_125_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_37_io_to_pes_4_out_bits = PE_125_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_37_io_to_pes_4_in_ready = PE_125_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_37_io_to_pes_5_out_valid = PE_126_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_37_io_to_pes_5_out_bits = PE_126_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_37_io_to_pes_5_in_ready = PE_126_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_37_io_to_pes_6_out_valid = PE_127_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_37_io_to_pes_6_out_bits = PE_127_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_37_io_to_pes_6_in_ready = PE_127_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_37_io_to_pes_7_out_valid = PE_128_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_37_io_to_pes_7_out_bits = PE_128_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_37_io_to_pes_7_in_ready = PE_128_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_37_io_to_pes_8_out_valid = PE_129_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_37_io_to_pes_8_out_bits = PE_129_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_37_io_to_pes_8_in_ready = PE_129_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_37_io_to_pes_9_out_valid = PE_130_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_37_io_to_pes_9_out_bits = PE_130_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_37_io_to_pes_9_in_ready = PE_130_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_37_io_to_pes_10_out_valid = PE_131_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_37_io_to_pes_10_out_bits = PE_131_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_37_io_to_pes_10_in_ready = PE_131_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_37_io_sig_stat2trans = MultiDimTime_io_index_1 == 16'h0; // @[pe.scala 281:43]
  assign PENetwork_38_clock = clock;
  assign PENetwork_38_io_to_pes_0_out_valid = PE_132_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_38_io_to_pes_0_out_bits = PE_132_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_38_io_to_pes_1_out_valid = PE_133_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_38_io_to_pes_1_out_bits = PE_133_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_38_io_to_pes_1_in_ready = PE_133_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_38_io_to_pes_2_out_valid = PE_134_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_38_io_to_pes_2_out_bits = PE_134_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_38_io_to_pes_2_in_ready = PE_134_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_38_io_to_pes_3_out_valid = PE_135_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_38_io_to_pes_3_out_bits = PE_135_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_38_io_to_pes_3_in_ready = PE_135_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_38_io_to_pes_4_out_valid = PE_136_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_38_io_to_pes_4_out_bits = PE_136_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_38_io_to_pes_4_in_ready = PE_136_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_38_io_to_pes_5_out_valid = PE_137_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_38_io_to_pes_5_out_bits = PE_137_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_38_io_to_pes_5_in_ready = PE_137_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_38_io_to_pes_6_out_valid = PE_138_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_38_io_to_pes_6_out_bits = PE_138_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_38_io_to_pes_6_in_ready = PE_138_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_38_io_to_pes_7_out_valid = PE_139_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_38_io_to_pes_7_out_bits = PE_139_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_38_io_to_pes_7_in_ready = PE_139_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_38_io_to_pes_8_out_valid = PE_140_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_38_io_to_pes_8_out_bits = PE_140_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_38_io_to_pes_8_in_ready = PE_140_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_38_io_to_pes_9_out_valid = PE_141_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_38_io_to_pes_9_out_bits = PE_141_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_38_io_to_pes_9_in_ready = PE_141_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_38_io_to_pes_10_out_valid = PE_142_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_38_io_to_pes_10_out_bits = PE_142_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_38_io_to_pes_10_in_ready = PE_142_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_38_io_sig_stat2trans = MultiDimTime_io_index_1 == 16'h0; // @[pe.scala 281:43]
  assign PENetwork_39_clock = clock;
  assign PENetwork_39_io_to_pes_0_out_valid = PE_143_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_39_io_to_pes_0_out_bits = PE_143_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_39_io_to_pes_1_out_valid = PE_144_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_39_io_to_pes_1_out_bits = PE_144_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_39_io_to_pes_1_in_ready = PE_144_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_39_io_to_pes_2_out_valid = PE_145_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_39_io_to_pes_2_out_bits = PE_145_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_39_io_to_pes_2_in_ready = PE_145_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_39_io_to_pes_3_out_valid = PE_146_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_39_io_to_pes_3_out_bits = PE_146_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_39_io_to_pes_3_in_ready = PE_146_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_39_io_to_pes_4_out_valid = PE_147_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_39_io_to_pes_4_out_bits = PE_147_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_39_io_to_pes_4_in_ready = PE_147_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_39_io_to_pes_5_out_valid = PE_148_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_39_io_to_pes_5_out_bits = PE_148_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_39_io_to_pes_5_in_ready = PE_148_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_39_io_to_pes_6_out_valid = PE_149_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_39_io_to_pes_6_out_bits = PE_149_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_39_io_to_pes_6_in_ready = PE_149_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_39_io_to_pes_7_out_valid = PE_150_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_39_io_to_pes_7_out_bits = PE_150_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_39_io_to_pes_7_in_ready = PE_150_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_39_io_to_pes_8_out_valid = PE_151_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_39_io_to_pes_8_out_bits = PE_151_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_39_io_to_pes_8_in_ready = PE_151_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_39_io_to_pes_9_out_valid = PE_152_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_39_io_to_pes_9_out_bits = PE_152_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_39_io_to_pes_9_in_ready = PE_152_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_39_io_to_pes_10_out_valid = PE_153_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_39_io_to_pes_10_out_bits = PE_153_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_39_io_to_pes_10_in_ready = PE_153_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_39_io_sig_stat2trans = MultiDimTime_io_index_1 == 16'h0; // @[pe.scala 281:43]
  assign PENetwork_40_clock = clock;
  assign PENetwork_40_io_to_pes_0_out_valid = PE_154_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_40_io_to_pes_0_out_bits = PE_154_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_40_io_to_pes_1_out_valid = PE_155_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_40_io_to_pes_1_out_bits = PE_155_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_40_io_to_pes_1_in_ready = PE_155_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_40_io_to_pes_2_out_valid = PE_156_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_40_io_to_pes_2_out_bits = PE_156_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_40_io_to_pes_2_in_ready = PE_156_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_40_io_to_pes_3_out_valid = PE_157_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_40_io_to_pes_3_out_bits = PE_157_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_40_io_to_pes_3_in_ready = PE_157_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_40_io_to_pes_4_out_valid = PE_158_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_40_io_to_pes_4_out_bits = PE_158_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_40_io_to_pes_4_in_ready = PE_158_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_40_io_to_pes_5_out_valid = PE_159_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_40_io_to_pes_5_out_bits = PE_159_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_40_io_to_pes_5_in_ready = PE_159_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_40_io_to_pes_6_out_valid = PE_160_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_40_io_to_pes_6_out_bits = PE_160_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_40_io_to_pes_6_in_ready = PE_160_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_40_io_to_pes_7_out_valid = PE_161_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_40_io_to_pes_7_out_bits = PE_161_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_40_io_to_pes_7_in_ready = PE_161_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_40_io_to_pes_8_out_valid = PE_162_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_40_io_to_pes_8_out_bits = PE_162_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_40_io_to_pes_8_in_ready = PE_162_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_40_io_to_pes_9_out_valid = PE_163_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_40_io_to_pes_9_out_bits = PE_163_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_40_io_to_pes_9_in_ready = PE_163_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_40_io_to_pes_10_out_valid = PE_164_io_data_2_out_valid; // @[pe.scala 261:36]
  assign PENetwork_40_io_to_pes_10_out_bits = PE_164_io_data_2_out_bits; // @[pe.scala 261:36]
  assign PENetwork_40_io_to_pes_10_in_ready = PE_164_io_data_2_in_ready; // @[pe.scala 267:49]
  assign PENetwork_40_io_sig_stat2trans = MultiDimTime_io_index_1 == 16'h0; // @[pe.scala 281:43]
  assign MemController_clock = clock;
  assign MemController_reset = reset;
  assign MemController_io_rd_valid = io_exec_valid; // @[pe.scala 313:28]
  assign MemController_io_wr_valid = io_data_0_in_0_valid; // @[pe.scala 314:28]
  assign MemController_io_wr_data_valid = io_data_0_in_0_bits_valid; // @[pe.scala 316:27]
  assign MemController_io_wr_data_bits = io_data_0_in_0_bits_bits; // @[pe.scala 316:27]
  assign MemController_1_clock = clock;
  assign MemController_1_reset = reset;
  assign MemController_1_io_rd_valid = io_exec_valid; // @[pe.scala 313:28]
  assign MemController_1_io_wr_valid = io_data_0_in_1_valid; // @[pe.scala 314:28]
  assign MemController_1_io_wr_data_valid = io_data_0_in_1_bits_valid; // @[pe.scala 316:27]
  assign MemController_1_io_wr_data_bits = io_data_0_in_1_bits_bits; // @[pe.scala 316:27]
  assign MemController_2_clock = clock;
  assign MemController_2_reset = reset;
  assign MemController_2_io_rd_valid = io_exec_valid; // @[pe.scala 313:28]
  assign MemController_2_io_wr_valid = io_data_0_in_2_valid; // @[pe.scala 314:28]
  assign MemController_2_io_wr_data_valid = io_data_0_in_2_bits_valid; // @[pe.scala 316:27]
  assign MemController_2_io_wr_data_bits = io_data_0_in_2_bits_bits; // @[pe.scala 316:27]
  assign MemController_3_clock = clock;
  assign MemController_3_reset = reset;
  assign MemController_3_io_rd_valid = io_exec_valid; // @[pe.scala 313:28]
  assign MemController_3_io_wr_valid = io_data_0_in_3_valid; // @[pe.scala 314:28]
  assign MemController_3_io_wr_data_valid = io_data_0_in_3_bits_valid; // @[pe.scala 316:27]
  assign MemController_3_io_wr_data_bits = io_data_0_in_3_bits_bits; // @[pe.scala 316:27]
  assign MemController_4_clock = clock;
  assign MemController_4_reset = reset;
  assign MemController_4_io_rd_valid = io_exec_valid; // @[pe.scala 313:28]
  assign MemController_4_io_wr_valid = io_data_0_in_4_valid; // @[pe.scala 314:28]
  assign MemController_4_io_wr_data_valid = io_data_0_in_4_bits_valid; // @[pe.scala 316:27]
  assign MemController_4_io_wr_data_bits = io_data_0_in_4_bits_bits; // @[pe.scala 316:27]
  assign MemController_5_clock = clock;
  assign MemController_5_reset = reset;
  assign MemController_5_io_rd_valid = io_exec_valid; // @[pe.scala 313:28]
  assign MemController_5_io_wr_valid = io_data_0_in_5_valid; // @[pe.scala 314:28]
  assign MemController_5_io_wr_data_valid = io_data_0_in_5_bits_valid; // @[pe.scala 316:27]
  assign MemController_5_io_wr_data_bits = io_data_0_in_5_bits_bits; // @[pe.scala 316:27]
  assign MemController_6_clock = clock;
  assign MemController_6_reset = reset;
  assign MemController_6_io_rd_valid = io_exec_valid; // @[pe.scala 313:28]
  assign MemController_6_io_wr_valid = io_data_0_in_6_valid; // @[pe.scala 314:28]
  assign MemController_6_io_wr_data_valid = io_data_0_in_6_bits_valid; // @[pe.scala 316:27]
  assign MemController_6_io_wr_data_bits = io_data_0_in_6_bits_bits; // @[pe.scala 316:27]
  assign MemController_7_clock = clock;
  assign MemController_7_reset = reset;
  assign MemController_7_io_rd_valid = io_exec_valid; // @[pe.scala 313:28]
  assign MemController_7_io_wr_valid = io_data_0_in_7_valid; // @[pe.scala 314:28]
  assign MemController_7_io_wr_data_valid = io_data_0_in_7_bits_valid; // @[pe.scala 316:27]
  assign MemController_7_io_wr_data_bits = io_data_0_in_7_bits_bits; // @[pe.scala 316:27]
  assign MemController_8_clock = clock;
  assign MemController_8_reset = reset;
  assign MemController_8_io_rd_valid = io_exec_valid; // @[pe.scala 313:28]
  assign MemController_8_io_wr_valid = io_data_0_in_8_valid; // @[pe.scala 314:28]
  assign MemController_8_io_wr_data_valid = io_data_0_in_8_bits_valid; // @[pe.scala 316:27]
  assign MemController_8_io_wr_data_bits = io_data_0_in_8_bits_bits; // @[pe.scala 316:27]
  assign MemController_9_clock = clock;
  assign MemController_9_reset = reset;
  assign MemController_9_io_rd_valid = io_exec_valid; // @[pe.scala 313:28]
  assign MemController_9_io_wr_valid = io_data_0_in_9_valid; // @[pe.scala 314:28]
  assign MemController_9_io_wr_data_valid = io_data_0_in_9_bits_valid; // @[pe.scala 316:27]
  assign MemController_9_io_wr_data_bits = io_data_0_in_9_bits_bits; // @[pe.scala 316:27]
  assign MemController_10_clock = clock;
  assign MemController_10_reset = reset;
  assign MemController_10_io_rd_valid = io_exec_valid; // @[pe.scala 313:28]
  assign MemController_10_io_wr_valid = io_data_0_in_10_valid; // @[pe.scala 314:28]
  assign MemController_10_io_wr_data_valid = io_data_0_in_10_bits_valid; // @[pe.scala 316:27]
  assign MemController_10_io_wr_data_bits = io_data_0_in_10_bits_bits; // @[pe.scala 316:27]
  assign MemController_11_clock = clock;
  assign MemController_11_reset = reset;
  assign MemController_11_io_rd_valid = io_exec_valid; // @[pe.scala 313:28]
  assign MemController_11_io_wr_valid = io_data_1_in_0_valid; // @[pe.scala 314:28]
  assign MemController_11_io_wr_data_valid = io_data_1_in_0_bits_valid; // @[pe.scala 316:27]
  assign MemController_11_io_wr_data_bits = io_data_1_in_0_bits_bits; // @[pe.scala 316:27]
  assign MemController_12_clock = clock;
  assign MemController_12_reset = reset;
  assign MemController_12_io_rd_valid = io_exec_valid; // @[pe.scala 313:28]
  assign MemController_12_io_wr_valid = io_data_1_in_1_valid; // @[pe.scala 314:28]
  assign MemController_12_io_wr_data_valid = io_data_1_in_1_bits_valid; // @[pe.scala 316:27]
  assign MemController_12_io_wr_data_bits = io_data_1_in_1_bits_bits; // @[pe.scala 316:27]
  assign MemController_13_clock = clock;
  assign MemController_13_reset = reset;
  assign MemController_13_io_rd_valid = io_exec_valid; // @[pe.scala 313:28]
  assign MemController_13_io_wr_valid = io_data_1_in_2_valid; // @[pe.scala 314:28]
  assign MemController_13_io_wr_data_valid = io_data_1_in_2_bits_valid; // @[pe.scala 316:27]
  assign MemController_13_io_wr_data_bits = io_data_1_in_2_bits_bits; // @[pe.scala 316:27]
  assign MemController_14_clock = clock;
  assign MemController_14_reset = reset;
  assign MemController_14_io_rd_valid = io_exec_valid; // @[pe.scala 313:28]
  assign MemController_14_io_wr_valid = io_data_1_in_3_valid; // @[pe.scala 314:28]
  assign MemController_14_io_wr_data_valid = io_data_1_in_3_bits_valid; // @[pe.scala 316:27]
  assign MemController_14_io_wr_data_bits = io_data_1_in_3_bits_bits; // @[pe.scala 316:27]
  assign MemController_15_clock = clock;
  assign MemController_15_reset = reset;
  assign MemController_15_io_rd_valid = io_exec_valid; // @[pe.scala 313:28]
  assign MemController_15_io_wr_valid = io_data_1_in_4_valid; // @[pe.scala 314:28]
  assign MemController_15_io_wr_data_valid = io_data_1_in_4_bits_valid; // @[pe.scala 316:27]
  assign MemController_15_io_wr_data_bits = io_data_1_in_4_bits_bits; // @[pe.scala 316:27]
  assign MemController_16_clock = clock;
  assign MemController_16_reset = reset;
  assign MemController_16_io_rd_valid = io_exec_valid; // @[pe.scala 313:28]
  assign MemController_16_io_wr_valid = io_data_1_in_5_valid; // @[pe.scala 314:28]
  assign MemController_16_io_wr_data_valid = io_data_1_in_5_bits_valid; // @[pe.scala 316:27]
  assign MemController_16_io_wr_data_bits = io_data_1_in_5_bits_bits; // @[pe.scala 316:27]
  assign MemController_17_clock = clock;
  assign MemController_17_reset = reset;
  assign MemController_17_io_rd_valid = io_exec_valid; // @[pe.scala 313:28]
  assign MemController_17_io_wr_valid = io_data_1_in_6_valid; // @[pe.scala 314:28]
  assign MemController_17_io_wr_data_valid = io_data_1_in_6_bits_valid; // @[pe.scala 316:27]
  assign MemController_17_io_wr_data_bits = io_data_1_in_6_bits_bits; // @[pe.scala 316:27]
  assign MemController_18_clock = clock;
  assign MemController_18_reset = reset;
  assign MemController_18_io_rd_valid = io_exec_valid; // @[pe.scala 313:28]
  assign MemController_18_io_wr_valid = io_data_1_in_7_valid; // @[pe.scala 314:28]
  assign MemController_18_io_wr_data_valid = io_data_1_in_7_bits_valid; // @[pe.scala 316:27]
  assign MemController_18_io_wr_data_bits = io_data_1_in_7_bits_bits; // @[pe.scala 316:27]
  assign MemController_19_clock = clock;
  assign MemController_19_reset = reset;
  assign MemController_19_io_rd_valid = io_exec_valid; // @[pe.scala 313:28]
  assign MemController_19_io_wr_valid = io_data_1_in_8_valid; // @[pe.scala 314:28]
  assign MemController_19_io_wr_data_valid = io_data_1_in_8_bits_valid; // @[pe.scala 316:27]
  assign MemController_19_io_wr_data_bits = io_data_1_in_8_bits_bits; // @[pe.scala 316:27]
  assign MemController_20_clock = clock;
  assign MemController_20_reset = reset;
  assign MemController_20_io_rd_valid = io_exec_valid; // @[pe.scala 313:28]
  assign MemController_20_io_wr_valid = io_data_1_in_9_valid; // @[pe.scala 314:28]
  assign MemController_20_io_wr_data_valid = io_data_1_in_9_bits_valid; // @[pe.scala 316:27]
  assign MemController_20_io_wr_data_bits = io_data_1_in_9_bits_bits; // @[pe.scala 316:27]
  assign MemController_21_clock = clock;
  assign MemController_21_reset = reset;
  assign MemController_21_io_rd_valid = io_exec_valid; // @[pe.scala 313:28]
  assign MemController_21_io_wr_valid = io_data_1_in_10_valid; // @[pe.scala 314:28]
  assign MemController_21_io_wr_data_valid = io_data_1_in_10_bits_valid; // @[pe.scala 316:27]
  assign MemController_21_io_wr_data_bits = io_data_1_in_10_bits_bits; // @[pe.scala 316:27]
  assign MemController_22_clock = clock;
  assign MemController_22_reset = reset;
  assign MemController_22_io_rd_valid = io_exec_valid; // @[pe.scala 313:28]
  assign MemController_22_io_wr_valid = io_data_1_in_11_valid; // @[pe.scala 314:28]
  assign MemController_22_io_wr_data_valid = io_data_1_in_11_bits_valid; // @[pe.scala 316:27]
  assign MemController_22_io_wr_data_bits = io_data_1_in_11_bits_bits; // @[pe.scala 316:27]
  assign MemController_23_clock = clock;
  assign MemController_23_reset = reset;
  assign MemController_23_io_rd_valid = io_exec_valid; // @[pe.scala 313:28]
  assign MemController_23_io_wr_valid = io_data_1_in_12_valid; // @[pe.scala 314:28]
  assign MemController_23_io_wr_data_valid = io_data_1_in_12_bits_valid; // @[pe.scala 316:27]
  assign MemController_23_io_wr_data_bits = io_data_1_in_12_bits_bits; // @[pe.scala 316:27]
  assign MemController_24_clock = clock;
  assign MemController_24_reset = reset;
  assign MemController_24_io_rd_valid = io_exec_valid; // @[pe.scala 313:28]
  assign MemController_24_io_wr_valid = io_data_1_in_13_valid; // @[pe.scala 314:28]
  assign MemController_24_io_wr_data_valid = io_data_1_in_13_bits_valid; // @[pe.scala 316:27]
  assign MemController_24_io_wr_data_bits = io_data_1_in_13_bits_bits; // @[pe.scala 316:27]
  assign MemController_25_clock = clock;
  assign MemController_25_reset = reset;
  assign MemController_25_io_rd_valid = io_exec_valid; // @[pe.scala 313:28]
  assign MemController_25_io_wr_valid = io_data_1_in_14_valid; // @[pe.scala 314:28]
  assign MemController_25_io_wr_data_valid = io_data_1_in_14_bits_valid; // @[pe.scala 316:27]
  assign MemController_25_io_wr_data_bits = io_data_1_in_14_bits_bits; // @[pe.scala 316:27]
  assign MemController_26_clock = clock;
  assign MemController_26_reset = reset;
  assign MemController_26_io_rd_valid = io_out_valid; // @[pe.scala 319:28]
  assign MemController_26_io_wr_valid = PENetwork_26_io_to_mem_valid; // @[pe.scala 318:28]
  assign MemController_26_io_wr_data_valid = PENetwork_26_io_to_mem_valid; // @[pe.scala 320:27]
  assign MemController_26_io_wr_data_bits = PENetwork_26_io_to_mem_bits; // @[pe.scala 320:27]
  assign MemController_27_clock = clock;
  assign MemController_27_reset = reset;
  assign MemController_27_io_rd_valid = io_out_valid; // @[pe.scala 319:28]
  assign MemController_27_io_wr_valid = PENetwork_27_io_to_mem_valid; // @[pe.scala 318:28]
  assign MemController_27_io_wr_data_valid = PENetwork_27_io_to_mem_valid; // @[pe.scala 320:27]
  assign MemController_27_io_wr_data_bits = PENetwork_27_io_to_mem_bits; // @[pe.scala 320:27]
  assign MemController_28_clock = clock;
  assign MemController_28_reset = reset;
  assign MemController_28_io_rd_valid = io_out_valid; // @[pe.scala 319:28]
  assign MemController_28_io_wr_valid = PENetwork_28_io_to_mem_valid; // @[pe.scala 318:28]
  assign MemController_28_io_wr_data_valid = PENetwork_28_io_to_mem_valid; // @[pe.scala 320:27]
  assign MemController_28_io_wr_data_bits = PENetwork_28_io_to_mem_bits; // @[pe.scala 320:27]
  assign MemController_29_clock = clock;
  assign MemController_29_reset = reset;
  assign MemController_29_io_rd_valid = io_out_valid; // @[pe.scala 319:28]
  assign MemController_29_io_wr_valid = PENetwork_29_io_to_mem_valid; // @[pe.scala 318:28]
  assign MemController_29_io_wr_data_valid = PENetwork_29_io_to_mem_valid; // @[pe.scala 320:27]
  assign MemController_29_io_wr_data_bits = PENetwork_29_io_to_mem_bits; // @[pe.scala 320:27]
  assign MemController_30_clock = clock;
  assign MemController_30_reset = reset;
  assign MemController_30_io_rd_valid = io_out_valid; // @[pe.scala 319:28]
  assign MemController_30_io_wr_valid = PENetwork_30_io_to_mem_valid; // @[pe.scala 318:28]
  assign MemController_30_io_wr_data_valid = PENetwork_30_io_to_mem_valid; // @[pe.scala 320:27]
  assign MemController_30_io_wr_data_bits = PENetwork_30_io_to_mem_bits; // @[pe.scala 320:27]
  assign MemController_31_clock = clock;
  assign MemController_31_reset = reset;
  assign MemController_31_io_rd_valid = io_out_valid; // @[pe.scala 319:28]
  assign MemController_31_io_wr_valid = PENetwork_31_io_to_mem_valid; // @[pe.scala 318:28]
  assign MemController_31_io_wr_data_valid = PENetwork_31_io_to_mem_valid; // @[pe.scala 320:27]
  assign MemController_31_io_wr_data_bits = PENetwork_31_io_to_mem_bits; // @[pe.scala 320:27]
  assign MemController_32_clock = clock;
  assign MemController_32_reset = reset;
  assign MemController_32_io_rd_valid = io_out_valid; // @[pe.scala 319:28]
  assign MemController_32_io_wr_valid = PENetwork_32_io_to_mem_valid; // @[pe.scala 318:28]
  assign MemController_32_io_wr_data_valid = PENetwork_32_io_to_mem_valid; // @[pe.scala 320:27]
  assign MemController_32_io_wr_data_bits = PENetwork_32_io_to_mem_bits; // @[pe.scala 320:27]
  assign MemController_33_clock = clock;
  assign MemController_33_reset = reset;
  assign MemController_33_io_rd_valid = io_out_valid; // @[pe.scala 319:28]
  assign MemController_33_io_wr_valid = PENetwork_33_io_to_mem_valid; // @[pe.scala 318:28]
  assign MemController_33_io_wr_data_valid = PENetwork_33_io_to_mem_valid; // @[pe.scala 320:27]
  assign MemController_33_io_wr_data_bits = PENetwork_33_io_to_mem_bits; // @[pe.scala 320:27]
  assign MemController_34_clock = clock;
  assign MemController_34_reset = reset;
  assign MemController_34_io_rd_valid = io_out_valid; // @[pe.scala 319:28]
  assign MemController_34_io_wr_valid = PENetwork_34_io_to_mem_valid; // @[pe.scala 318:28]
  assign MemController_34_io_wr_data_valid = PENetwork_34_io_to_mem_valid; // @[pe.scala 320:27]
  assign MemController_34_io_wr_data_bits = PENetwork_34_io_to_mem_bits; // @[pe.scala 320:27]
  assign MemController_35_clock = clock;
  assign MemController_35_reset = reset;
  assign MemController_35_io_rd_valid = io_out_valid; // @[pe.scala 319:28]
  assign MemController_35_io_wr_valid = PENetwork_35_io_to_mem_valid; // @[pe.scala 318:28]
  assign MemController_35_io_wr_data_valid = PENetwork_35_io_to_mem_valid; // @[pe.scala 320:27]
  assign MemController_35_io_wr_data_bits = PENetwork_35_io_to_mem_bits; // @[pe.scala 320:27]
  assign MemController_36_clock = clock;
  assign MemController_36_reset = reset;
  assign MemController_36_io_rd_valid = io_out_valid; // @[pe.scala 319:28]
  assign MemController_36_io_wr_valid = PENetwork_36_io_to_mem_valid; // @[pe.scala 318:28]
  assign MemController_36_io_wr_data_valid = PENetwork_36_io_to_mem_valid; // @[pe.scala 320:27]
  assign MemController_36_io_wr_data_bits = PENetwork_36_io_to_mem_bits; // @[pe.scala 320:27]
  assign MemController_37_clock = clock;
  assign MemController_37_reset = reset;
  assign MemController_37_io_rd_valid = io_out_valid; // @[pe.scala 319:28]
  assign MemController_37_io_wr_valid = PENetwork_37_io_to_mem_valid; // @[pe.scala 318:28]
  assign MemController_37_io_wr_data_valid = PENetwork_37_io_to_mem_valid; // @[pe.scala 320:27]
  assign MemController_37_io_wr_data_bits = PENetwork_37_io_to_mem_bits; // @[pe.scala 320:27]
  assign MemController_38_clock = clock;
  assign MemController_38_reset = reset;
  assign MemController_38_io_rd_valid = io_out_valid; // @[pe.scala 319:28]
  assign MemController_38_io_wr_valid = PENetwork_38_io_to_mem_valid; // @[pe.scala 318:28]
  assign MemController_38_io_wr_data_valid = PENetwork_38_io_to_mem_valid; // @[pe.scala 320:27]
  assign MemController_38_io_wr_data_bits = PENetwork_38_io_to_mem_bits; // @[pe.scala 320:27]
  assign MemController_39_clock = clock;
  assign MemController_39_reset = reset;
  assign MemController_39_io_rd_valid = io_out_valid; // @[pe.scala 319:28]
  assign MemController_39_io_wr_valid = PENetwork_39_io_to_mem_valid; // @[pe.scala 318:28]
  assign MemController_39_io_wr_data_valid = PENetwork_39_io_to_mem_valid; // @[pe.scala 320:27]
  assign MemController_39_io_wr_data_bits = PENetwork_39_io_to_mem_bits; // @[pe.scala 320:27]
  assign MemController_40_clock = clock;
  assign MemController_40_reset = reset;
  assign MemController_40_io_rd_valid = io_out_valid; // @[pe.scala 319:28]
  assign MemController_40_io_wr_valid = PENetwork_40_io_to_mem_valid; // @[pe.scala 318:28]
  assign MemController_40_io_wr_data_valid = PENetwork_40_io_to_mem_valid; // @[pe.scala 320:27]
  assign MemController_40_io_wr_data_bits = PENetwork_40_io_to_mem_bits; // @[pe.scala 320:27]
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1) begin
          $fwrite(32'h80000002,"time_ctrl: %d %d %d\n",MultiDimTime_io_index_0,MultiDimTime_io_index_1,MultiDimTime_io_index_2); // @[pe.scala 163:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
