module MultiDimTime(
  input         clock,
  input         reset,
  input         io_in,
  output [1:0]  io_out_0,
  output [1:0]  io_out_1,
  output [17:0] io_index_0,
  output [17:0] io_index_1
);
  reg [15:0] regs_0; // @[mem.scala 67:12]
  reg [31:0] _RAND_0;
  reg [15:0] regs_1; // @[mem.scala 67:12]
  reg [31:0] _RAND_1;
  wire [15:0] _GEN_4 = {{15'd0}, io_in}; // @[mem.scala 69:42]
  wire [15:0] _T_1 = regs_0 + _GEN_4; // @[mem.scala 69:42]
  wire  back_0 = _T_1 == 16'h1; // @[mem.scala 69:48]
  wire [15:0] _T_3 = regs_1 + _GEN_4; // @[mem.scala 69:42]
  wire  back_1 = _T_3 == 16'h8; // @[mem.scala 69:48]
  wire  _T_4 = ~back_0; // @[mem.scala 76:20]
  wire [1:0] _T_5 = {_T_4, 1'h0}; // @[mem.scala 76:31]
  wire  _T_6 = ~back_1; // @[mem.scala 76:40]
  wire [1:0] _GEN_6 = {{1'd0}, _T_6}; // @[mem.scala 76:37]
  wire  _GEN_3 = back_0 ? 1'h0 : io_in; // @[mem.scala 86:16]
  assign io_out_0 = {{1'd0}, _GEN_3}; // @[mem.scala 88:15 mem.scala 91:15]
  assign io_out_1 = _T_5 | _GEN_6; // @[mem.scala 76:15]
  assign io_index_0 = {{2'd0}, regs_0}; // @[mem.scala 85:15]
  assign io_index_1 = {{2'd0}, regs_1}; // @[mem.scala 73:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 16'h0;
    end else if (back_0) begin
      regs_0 <= 16'h0;
    end else begin
      regs_0 <= _T_1;
    end
    if (reset) begin
      regs_1 <= 16'h0;
    end else if (back_0) begin
      if (back_1) begin
        regs_1 <= 16'h0;
      end else begin
        regs_1 <= _T_3;
      end
    end
  end
endmodule
module ComputeCell_Latency(
  input         clock,
  input         reset,
  input  [15:0] io_data_2_in,
  input  [15:0] io_data_1_in,
  input  [15:0] io_data_0_in,
  output [15:0] io_data_0_out
);
  reg [15:0] delay_a_0; // @[Reg.scala 27:20]
  reg [31:0] _RAND_0;
  reg [15:0] delay_b_0; // @[Reg.scala 27:20]
  reg [31:0] _RAND_1;
  reg [15:0] delay_c_0; // @[Reg.scala 27:20]
  reg [31:0] _RAND_2;
  wire [31:0] _T_9 = delay_a_0 * delay_b_0; // @[cell.scala 135:63]
  wire [31:0] _GEN_3 = {{16'd0}, delay_c_0}; // @[cell.scala 135:50]
  wire [31:0] _T_11 = _GEN_3 + _T_9; // @[cell.scala 135:50]
  assign io_data_0_out = _T_11[15:0]; // @[cell.scala 138:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  delay_a_0 = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  delay_b_0 = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  delay_c_0 = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      delay_a_0 <= 16'h0;
    end else begin
      delay_a_0 <= io_data_1_in;
    end
    if (reset) begin
      delay_b_0 <= 16'h0;
    end else begin
      delay_b_0 <= io_data_2_in;
    end
    if (reset) begin
      delay_c_0 <= 16'h0;
    end else begin
      delay_c_0 <= io_data_0_in;
    end
  end
endmodule
module SystolicOutput(
  input         io_port_in_valid,
  input  [15:0] io_port_in_bits,
  output        io_port_out_valid,
  output [15:0] io_port_out_bits,
  input         io_from_cell_valid,
  input  [15:0] io_from_cell_bits,
  output        io_to_cell_valid,
  output [15:0] io_to_cell_bits
);
  assign io_port_out_valid = io_from_cell_valid; // @[pe_modules.scala 111:15]
  assign io_port_out_bits = io_from_cell_bits; // @[pe_modules.scala 111:15]
  assign io_to_cell_valid = io_port_in_valid; // @[pe_modules.scala 110:14]
  assign io_to_cell_bits = io_port_in_bits; // @[pe_modules.scala 110:14]
endmodule
module StationaryInput_Pipeline(
  input         clock,
  input         reset,
  input         io_port_in_valid,
  input  [15:0] io_port_in_bits,
  output        io_port_out_valid,
  output [15:0] io_port_out_bits,
  output [15:0] io_to_cell_bits,
  input         io_sig_stat2trans
);
  reg  trans_valid; // @[pe_modules.scala 128:22]
  reg [31:0] _RAND_0;
  reg [15:0] trans_bits; // @[pe_modules.scala 128:22]
  reg [31:0] _RAND_1;
  reg  update_valid; // @[pe_modules.scala 131:23]
  reg [31:0] _RAND_2;
  reg [15:0] update_bits_0; // @[pe_modules.scala 131:23]
  reg [31:0] _RAND_3;
  reg [15:0] stat_bits_0; // @[pe_modules.scala 133:21]
  reg [31:0] _RAND_4;
  reg  reg_stat2trans_0; // @[pe_modules.scala 135:31]
  reg [31:0] _RAND_5;
  reg [3:0] write_trans_pos; // @[pe_modules.scala 137:32]
  reg [31:0] _RAND_6;
  wire  _T_4 = ~update_valid; // @[pe_modules.scala 142:26]
  wire [3:0] _GEN_5 = {{3'd0}, trans_valid}; // @[pe_modules.scala 142:60]
  wire [3:0] _T_6 = write_trans_pos + _GEN_5; // @[pe_modules.scala 142:60]
  wire  _T_7 = _T_6 == 4'h1; // @[pe_modules.scala 142:79]
  wire  _T_13 = _T_4 & trans_valid; // @[pe_modules.scala 143:24]
  wire  _T_21 = write_trans_pos == 4'h0; // @[pe_modules.scala 149:23]
  wire  _T_22 = _T_21 & trans_valid; // @[pe_modules.scala 149:45]
  wire  _GEN_1 = _T_22 | update_valid; // @[pe_modules.scala 149:60]
  reg [15:0] _T_24; // @[pe_modules.scala 163:29]
  reg [31:0] _RAND_7;
  assign io_port_out_valid = update_valid; // @[pe_modules.scala 139:21]
  assign io_port_out_bits = trans_bits; // @[pe_modules.scala 140:20]
  assign io_to_cell_bits = _T_24; // @[pe_modules.scala 163:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  trans_valid = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  trans_bits = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  update_valid = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  update_bits_0 = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  stat_bits_0 = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  reg_stat2trans_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  write_trans_pos = _RAND_6[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_24 = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      trans_valid <= 1'h0;
    end else begin
      trans_valid <= io_port_in_valid;
    end
    if (reset) begin
      trans_bits <= 16'h0;
    end else begin
      trans_bits <= io_port_in_bits;
    end
    if (reset) begin
      update_valid <= 1'h0;
    end else if (reg_stat2trans_0) begin
      update_valid <= 1'h0;
    end else begin
      update_valid <= _GEN_1;
    end
    if (reset) begin
      update_bits_0 <= 16'h0;
    end else if (_T_13) begin
      update_bits_0 <= trans_bits;
    end
    if (reset) begin
      stat_bits_0 <= 16'h0;
    end else if (reg_stat2trans_0) begin
      stat_bits_0 <= update_bits_0;
    end
    if (reset) begin
      reg_stat2trans_0 <= 1'h0;
    end else begin
      reg_stat2trans_0 <= io_sig_stat2trans;
    end
    if (reset) begin
      write_trans_pos <= 4'h0;
    end else if (_T_4) begin
      if (_T_7) begin
        write_trans_pos <= 4'h0;
      end else begin
        write_trans_pos <= _T_6;
      end
    end
    if (reset) begin
      _T_24 <= 16'h0;
    end else begin
      _T_24 <= stat_bits_0;
    end
  end
endmodule
module SystolicInput(
  input         clock,
  input         reset,
  input         io_port_in_valid,
  input  [15:0] io_port_in_bits,
  output        io_port_out_valid,
  output [15:0] io_port_out_bits,
  output [15:0] io_to_cell_bits
);
  reg  reg_0_valid; // @[pe_modules.scala 82:20]
  reg [31:0] _RAND_0;
  reg [15:0] reg_0_bits; // @[pe_modules.scala 82:20]
  reg [31:0] _RAND_1;
  reg [15:0] to_cell_delay1_bits; // @[pe_modules.scala 83:31]
  reg [31:0] _RAND_2;
  reg [15:0] to_cell_delay2_bits; // @[pe_modules.scala 84:31]
  reg [31:0] _RAND_3;
  assign io_port_out_valid = reg_0_valid; // @[pe_modules.scala 91:15]
  assign io_port_out_bits = reg_0_bits; // @[pe_modules.scala 91:15]
  assign io_to_cell_bits = to_cell_delay2_bits; // @[pe_modules.scala 92:14]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_0_valid = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  reg_0_bits = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  to_cell_delay1_bits = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  to_cell_delay2_bits = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      reg_0_valid <= 1'h0;
    end else begin
      reg_0_valid <= io_port_in_valid;
    end
    if (reset) begin
      reg_0_bits <= 16'h0;
    end else begin
      reg_0_bits <= io_port_in_bits;
    end
    if (reset) begin
      to_cell_delay1_bits <= 16'h0;
    end else begin
      to_cell_delay1_bits <= reg_0_bits;
    end
    if (reset) begin
      to_cell_delay2_bits <= 16'h0;
    end else begin
      to_cell_delay2_bits <= to_cell_delay1_bits;
    end
  end
endmodule
module PE(
  input         clock,
  input         reset,
  input         io_data_2_in_valid,
  input  [15:0] io_data_2_in_bits,
  output        io_data_2_out_valid,
  output [15:0] io_data_2_out_bits,
  input         io_data_1_in_valid,
  input  [15:0] io_data_1_in_bits,
  output        io_data_1_out_valid,
  output [15:0] io_data_1_out_bits,
  input         io_data_0_in_valid,
  input  [15:0] io_data_0_in_bits,
  output        io_data_0_out_valid,
  output [15:0] io_data_0_out_bits,
  input         io_sig_stat2trans
);
  wire  ComputeCell_Latency_clock; // @[pe.scala 37:18]
  wire  ComputeCell_Latency_reset; // @[pe.scala 37:18]
  wire [15:0] ComputeCell_Latency_io_data_2_in; // @[pe.scala 37:18]
  wire [15:0] ComputeCell_Latency_io_data_1_in; // @[pe.scala 37:18]
  wire [15:0] ComputeCell_Latency_io_data_0_in; // @[pe.scala 37:18]
  wire [15:0] ComputeCell_Latency_io_data_0_out; // @[pe.scala 37:18]
  wire  SystolicOutput_io_port_in_valid; // @[pe.scala 39:11]
  wire [15:0] SystolicOutput_io_port_in_bits; // @[pe.scala 39:11]
  wire  SystolicOutput_io_port_out_valid; // @[pe.scala 39:11]
  wire [15:0] SystolicOutput_io_port_out_bits; // @[pe.scala 39:11]
  wire  SystolicOutput_io_from_cell_valid; // @[pe.scala 39:11]
  wire [15:0] SystolicOutput_io_from_cell_bits; // @[pe.scala 39:11]
  wire  SystolicOutput_io_to_cell_valid; // @[pe.scala 39:11]
  wire [15:0] SystolicOutput_io_to_cell_bits; // @[pe.scala 39:11]
  wire  StationaryInput_Pipeline_clock; // @[pe.scala 39:11]
  wire  StationaryInput_Pipeline_reset; // @[pe.scala 39:11]
  wire  StationaryInput_Pipeline_io_port_in_valid; // @[pe.scala 39:11]
  wire [15:0] StationaryInput_Pipeline_io_port_in_bits; // @[pe.scala 39:11]
  wire  StationaryInput_Pipeline_io_port_out_valid; // @[pe.scala 39:11]
  wire [15:0] StationaryInput_Pipeline_io_port_out_bits; // @[pe.scala 39:11]
  wire [15:0] StationaryInput_Pipeline_io_to_cell_bits; // @[pe.scala 39:11]
  wire  StationaryInput_Pipeline_io_sig_stat2trans; // @[pe.scala 39:11]
  wire  SystolicInput_clock; // @[pe.scala 39:11]
  wire  SystolicInput_reset; // @[pe.scala 39:11]
  wire  SystolicInput_io_port_in_valid; // @[pe.scala 39:11]
  wire [15:0] SystolicInput_io_port_in_bits; // @[pe.scala 39:11]
  wire  SystolicInput_io_port_out_valid; // @[pe.scala 39:11]
  wire [15:0] SystolicInput_io_port_out_bits; // @[pe.scala 39:11]
  wire [15:0] SystolicInput_io_to_cell_bits; // @[pe.scala 39:11]
  reg  _T_3; // @[Reg.scala 15:16]
  reg [31:0] _RAND_0;
  ComputeCell_Latency ComputeCell_Latency ( // @[pe.scala 37:18]
    .clock(ComputeCell_Latency_clock),
    .reset(ComputeCell_Latency_reset),
    .io_data_2_in(ComputeCell_Latency_io_data_2_in),
    .io_data_1_in(ComputeCell_Latency_io_data_1_in),
    .io_data_0_in(ComputeCell_Latency_io_data_0_in),
    .io_data_0_out(ComputeCell_Latency_io_data_0_out)
  );
  SystolicOutput SystolicOutput ( // @[pe.scala 39:11]
    .io_port_in_valid(SystolicOutput_io_port_in_valid),
    .io_port_in_bits(SystolicOutput_io_port_in_bits),
    .io_port_out_valid(SystolicOutput_io_port_out_valid),
    .io_port_out_bits(SystolicOutput_io_port_out_bits),
    .io_from_cell_valid(SystolicOutput_io_from_cell_valid),
    .io_from_cell_bits(SystolicOutput_io_from_cell_bits),
    .io_to_cell_valid(SystolicOutput_io_to_cell_valid),
    .io_to_cell_bits(SystolicOutput_io_to_cell_bits)
  );
  StationaryInput_Pipeline StationaryInput_Pipeline ( // @[pe.scala 39:11]
    .clock(StationaryInput_Pipeline_clock),
    .reset(StationaryInput_Pipeline_reset),
    .io_port_in_valid(StationaryInput_Pipeline_io_port_in_valid),
    .io_port_in_bits(StationaryInput_Pipeline_io_port_in_bits),
    .io_port_out_valid(StationaryInput_Pipeline_io_port_out_valid),
    .io_port_out_bits(StationaryInput_Pipeline_io_port_out_bits),
    .io_to_cell_bits(StationaryInput_Pipeline_io_to_cell_bits),
    .io_sig_stat2trans(StationaryInput_Pipeline_io_sig_stat2trans)
  );
  SystolicInput SystolicInput ( // @[pe.scala 39:11]
    .clock(SystolicInput_clock),
    .reset(SystolicInput_reset),
    .io_port_in_valid(SystolicInput_io_port_in_valid),
    .io_port_in_bits(SystolicInput_io_port_in_bits),
    .io_port_out_valid(SystolicInput_io_port_out_valid),
    .io_port_out_bits(SystolicInput_io_port_out_bits),
    .io_to_cell_bits(SystolicInput_io_to_cell_bits)
  );
  assign io_data_2_out_valid = SystolicInput_io_port_out_valid; // @[pe.scala 42:17]
  assign io_data_2_out_bits = SystolicInput_io_port_out_bits; // @[pe.scala 42:17]
  assign io_data_1_out_valid = StationaryInput_Pipeline_io_port_out_valid; // @[pe.scala 42:17]
  assign io_data_1_out_bits = StationaryInput_Pipeline_io_port_out_bits; // @[pe.scala 42:17]
  assign io_data_0_out_valid = SystolicOutput_io_port_out_valid; // @[pe.scala 42:17]
  assign io_data_0_out_bits = SystolicOutput_io_port_out_bits; // @[pe.scala 42:17]
  assign ComputeCell_Latency_clock = clock;
  assign ComputeCell_Latency_reset = reset;
  assign ComputeCell_Latency_io_data_2_in = SystolicInput_io_to_cell_bits; // @[pe.scala 43:19]
  assign ComputeCell_Latency_io_data_1_in = StationaryInput_Pipeline_io_to_cell_bits; // @[pe.scala 43:19]
  assign ComputeCell_Latency_io_data_0_in = SystolicOutput_io_to_cell_bits; // @[pe.scala 43:19]
  assign SystolicOutput_io_port_in_valid = io_data_0_in_valid; // @[pe.scala 42:17]
  assign SystolicOutput_io_port_in_bits = io_data_0_in_bits; // @[pe.scala 42:17]
  assign SystolicOutput_io_from_cell_valid = _T_3; // @[pe.scala 46:34]
  assign SystolicOutput_io_from_cell_bits = ComputeCell_Latency_io_data_0_out; // @[pe.scala 45:33]
  assign StationaryInput_Pipeline_clock = clock;
  assign StationaryInput_Pipeline_reset = reset;
  assign StationaryInput_Pipeline_io_port_in_valid = io_data_1_in_valid; // @[pe.scala 42:17]
  assign StationaryInput_Pipeline_io_port_in_bits = io_data_1_in_bits; // @[pe.scala 42:17]
  assign StationaryInput_Pipeline_io_sig_stat2trans = io_sig_stat2trans; // @[pe.scala 50:33]
  assign SystolicInput_clock = clock;
  assign SystolicInput_reset = reset;
  assign SystolicInput_io_port_in_valid = io_data_2_in_valid; // @[pe.scala 42:17]
  assign SystolicInput_io_port_in_bits = io_data_2_in_bits; // @[pe.scala 42:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_3 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_3 <= SystolicOutput_io_to_cell_valid;
  end
endmodule
module PENetwork(
  input         io_to_pes_0_out_valid,
  input  [15:0] io_to_pes_0_out_bits,
  output        io_to_pes_1_in_valid,
  output [15:0] io_to_pes_1_in_bits,
  input         io_to_pes_1_out_valid,
  input  [15:0] io_to_pes_1_out_bits,
  output        io_to_pes_2_in_valid,
  output [15:0] io_to_pes_2_in_bits,
  input         io_to_pes_2_out_valid,
  input  [15:0] io_to_pes_2_out_bits,
  output        io_to_pes_3_in_valid,
  output [15:0] io_to_pes_3_in_bits,
  input         io_to_pes_3_out_valid,
  input  [15:0] io_to_pes_3_out_bits,
  output        io_to_pes_4_in_valid,
  output [15:0] io_to_pes_4_in_bits,
  input         io_to_pes_4_out_valid,
  input  [15:0] io_to_pes_4_out_bits,
  output        io_to_pes_5_in_valid,
  output [15:0] io_to_pes_5_in_bits,
  input         io_to_pes_5_out_valid,
  input  [15:0] io_to_pes_5_out_bits,
  output        io_to_pes_6_in_valid,
  output [15:0] io_to_pes_6_in_bits,
  input         io_to_pes_6_out_valid,
  input  [15:0] io_to_pes_6_out_bits,
  output        io_to_pes_7_in_valid,
  output [15:0] io_to_pes_7_in_bits,
  input         io_to_pes_7_out_valid,
  input  [15:0] io_to_pes_7_out_bits,
  output        io_to_mem_valid,
  output [15:0] io_to_mem_bits
);
  assign io_to_pes_1_in_valid = io_to_pes_0_out_valid; // @[pearray.scala 38:23]
  assign io_to_pes_1_in_bits = io_to_pes_0_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_2_in_valid = io_to_pes_1_out_valid; // @[pearray.scala 38:23]
  assign io_to_pes_2_in_bits = io_to_pes_1_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_3_in_valid = io_to_pes_2_out_valid; // @[pearray.scala 38:23]
  assign io_to_pes_3_in_bits = io_to_pes_2_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_4_in_valid = io_to_pes_3_out_valid; // @[pearray.scala 38:23]
  assign io_to_pes_4_in_bits = io_to_pes_3_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_5_in_valid = io_to_pes_4_out_valid; // @[pearray.scala 38:23]
  assign io_to_pes_5_in_bits = io_to_pes_4_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_6_in_valid = io_to_pes_5_out_valid; // @[pearray.scala 38:23]
  assign io_to_pes_6_in_bits = io_to_pes_5_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_7_in_valid = io_to_pes_6_out_valid; // @[pearray.scala 38:23]
  assign io_to_pes_7_in_bits = io_to_pes_6_out_bits; // @[pearray.scala 38:23]
  assign io_to_mem_valid = io_to_pes_7_out_valid; // @[pearray.scala 45:17]
  assign io_to_mem_bits = io_to_pes_7_out_bits; // @[pearray.scala 45:17]
endmodule
module PENetwork_8(
  output        io_to_pes_0_in_valid,
  output [15:0] io_to_pes_0_in_bits,
  input         io_to_pes_0_out_valid,
  input  [15:0] io_to_pes_0_out_bits,
  output        io_to_pes_1_in_valid,
  output [15:0] io_to_pes_1_in_bits,
  input         io_to_pes_1_out_valid,
  input  [15:0] io_to_pes_1_out_bits,
  output        io_to_pes_2_in_valid,
  output [15:0] io_to_pes_2_in_bits,
  input         io_to_pes_2_out_valid,
  input  [15:0] io_to_pes_2_out_bits,
  output        io_to_pes_3_in_valid,
  output [15:0] io_to_pes_3_in_bits,
  input         io_to_pes_3_out_valid,
  input  [15:0] io_to_pes_3_out_bits,
  output        io_to_pes_4_in_valid,
  output [15:0] io_to_pes_4_in_bits,
  input         io_to_pes_4_out_valid,
  input  [15:0] io_to_pes_4_out_bits,
  output        io_to_pes_5_in_valid,
  output [15:0] io_to_pes_5_in_bits,
  input         io_to_pes_5_out_valid,
  input  [15:0] io_to_pes_5_out_bits,
  output        io_to_pes_6_in_valid,
  output [15:0] io_to_pes_6_in_bits,
  input         io_to_pes_6_out_valid,
  input  [15:0] io_to_pes_6_out_bits,
  output        io_to_pes_7_in_valid,
  output [15:0] io_to_pes_7_in_bits,
  input         io_to_mem_valid,
  input  [15:0] io_to_mem_bits
);
  assign io_to_pes_0_in_valid = io_to_mem_valid; // @[pearray.scala 41:23]
  assign io_to_pes_0_in_bits = io_to_mem_bits; // @[pearray.scala 41:23]
  assign io_to_pes_1_in_valid = io_to_pes_0_out_valid; // @[pearray.scala 38:23]
  assign io_to_pes_1_in_bits = io_to_pes_0_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_2_in_valid = io_to_pes_1_out_valid; // @[pearray.scala 38:23]
  assign io_to_pes_2_in_bits = io_to_pes_1_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_3_in_valid = io_to_pes_2_out_valid; // @[pearray.scala 38:23]
  assign io_to_pes_3_in_bits = io_to_pes_2_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_4_in_valid = io_to_pes_3_out_valid; // @[pearray.scala 38:23]
  assign io_to_pes_4_in_bits = io_to_pes_3_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_5_in_valid = io_to_pes_4_out_valid; // @[pearray.scala 38:23]
  assign io_to_pes_5_in_bits = io_to_pes_4_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_6_in_valid = io_to_pes_5_out_valid; // @[pearray.scala 38:23]
  assign io_to_pes_6_in_bits = io_to_pes_5_out_bits; // @[pearray.scala 38:23]
  assign io_to_pes_7_in_valid = io_to_pes_6_out_valid; // @[pearray.scala 38:23]
  assign io_to_pes_7_in_bits = io_to_pes_6_out_bits; // @[pearray.scala 38:23]
endmodule
module MultiDimMem(
  input         clock,
  input         reset,
  input         io_rd_addr_valid,
  input  [1:0]  io_rd_addr_bits_0,
  input  [1:0]  io_rd_addr_bits_1,
  output        io_rd_data_valid,
  output [15:0] io_rd_data_bits,
  input  [1:0]  io_wr_addr_bits_0,
  input  [1:0]  io_wr_addr_bits_1,
  input         io_wr_data_valid,
  input  [15:0] io_wr_data_bits
);
  reg [16:0] mem [0:7]; // @[mem.scala 105:24]
  reg [31:0] _RAND_0;
  wire [16:0] mem_mem_output_data; // @[mem.scala 105:24]
  wire [2:0] mem_mem_output_addr; // @[mem.scala 105:24]
  wire [16:0] mem__T_43_data; // @[mem.scala 105:24]
  wire [2:0] mem__T_43_addr; // @[mem.scala 105:24]
  wire  mem__T_43_mask; // @[mem.scala 105:24]
  wire  mem__T_43_en; // @[mem.scala 105:24]
  reg  mem_mem_output_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [2:0] mem_mem_output_addr_pipe_0;
  reg [31:0] _RAND_2;
  reg  rd_addr_reg_valid; // @[mem.scala 106:28]
  reg [31:0] _RAND_3;
  reg [15:0] rd_addr_reg_bits_1; // @[mem.scala 106:28]
  reg [31:0] _RAND_4;
  reg [15:0] rd_addr_reg_bits_0; // @[mem.scala 106:28]
  reg [31:0] _RAND_5;
  wire [15:0] _T_6 = rd_addr_reg_bits_0 + 16'h1; // @[mem.scala 117:102]
  wire  _T_7 = 2'h1 == io_rd_addr_bits_0; // @[Mux.scala 68:19]
  wire  _T_9 = 2'h0 == io_rd_addr_bits_0; // @[Mux.scala 68:19]
  wire [15:0] _T_11 = rd_addr_reg_bits_1 + 16'h1; // @[mem.scala 117:102]
  wire  _T_12 = 2'h1 == io_rd_addr_bits_1; // @[Mux.scala 68:19]
  wire  _T_14 = 2'h0 == io_rd_addr_bits_1; // @[Mux.scala 68:19]
  wire [15:0] mem_rd_addr = rd_addr_reg_bits_0 + rd_addr_reg_bits_1; // @[mem.scala 120:46]
  reg  mem_req_valid; // @[mem.scala 125:30]
  reg [31:0] _RAND_6;
  reg [15:0] wr_addr_reg_bits_1; // @[mem.scala 126:28]
  reg [31:0] _RAND_7;
  reg [15:0] wr_addr_reg_bits_0; // @[mem.scala 126:28]
  reg [31:0] _RAND_8;
  wire [15:0] _T_22 = wr_addr_reg_bits_0 + 16'h1; // @[mem.scala 138:102]
  wire  _T_23 = 2'h1 == io_wr_addr_bits_0; // @[Mux.scala 68:19]
  wire  _T_25 = 2'h0 == io_wr_addr_bits_0; // @[Mux.scala 68:19]
  wire [15:0] _T_27 = wr_addr_reg_bits_1 + 16'h1; // @[mem.scala 138:102]
  wire  _T_28 = 2'h1 == io_wr_addr_bits_1; // @[Mux.scala 68:19]
  wire  _T_30 = 2'h0 == io_wr_addr_bits_1; // @[Mux.scala 68:19]
  wire [15:0] mem_wr_addr = wr_addr_reg_bits_0 + wr_addr_reg_bits_1; // @[mem.scala 140:46]
  reg  wr_data_1_valid; // @[mem.scala 145:26]
  reg [31:0] _RAND_9;
  reg [15:0] wr_data_1_bits; // @[mem.scala 145:26]
  reg [31:0] _RAND_10;
  reg  wr_data_2_valid; // @[mem.scala 152:26]
  reg [31:0] _RAND_11;
  reg [15:0] wr_data_2_bits; // @[mem.scala 152:26]
  reg [31:0] _RAND_12;
  reg [15:0] wr_addr_2; // @[mem.scala 154:26]
  reg [31:0] _RAND_13;
  reg [15:0] wr_data_final; // @[mem.scala 160:30]
  reg [31:0] _RAND_14;
  reg [15:0] wr_addr_3; // @[mem.scala 161:26]
  reg [31:0] _RAND_15;
  reg  wr_valid_3; // @[mem.scala 162:27]
  reg [31:0] _RAND_16;
  wire [16:0] _GEN_9 = {wr_valid_3, 16'h0}; // @[mem.scala 165:38]
  wire [31:0] _T_39 = {{15'd0}, _GEN_9}; // @[mem.scala 165:38]
  wire [31:0] _GEN_10 = {{16'd0}, wr_data_final}; // @[mem.scala 165:52]
  wire [31:0] _T_40 = _T_39 | _GEN_10; // @[mem.scala 165:52]
  reg  _T_46; // @[mem.scala 168:30]
  reg [31:0] _RAND_17;
  reg [15:0] _T_49; // @[mem.scala 169:29]
  reg [31:0] _RAND_18;
  assign mem_mem_output_addr = mem_mem_output_addr_pipe_0;
  assign mem_mem_output_data = mem[mem_mem_output_addr]; // @[mem.scala 105:24]
  assign mem__T_43_data = _T_40[16:0];
  assign mem__T_43_addr = wr_addr_3[2:0];
  assign mem__T_43_mask = 1'h1;
  assign mem__T_43_en = wr_valid_3;
  assign io_rd_data_valid = _T_46; // @[mem.scala 168:20]
  assign io_rd_data_bits = _T_49; // @[mem.scala 169:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    mem[initvar] = _RAND_0[16:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mem_mem_output_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  mem_mem_output_addr_pipe_0 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  rd_addr_reg_valid = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  rd_addr_reg_bits_1 = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  rd_addr_reg_bits_0 = _RAND_5[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  mem_req_valid = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  wr_addr_reg_bits_1 = _RAND_7[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  wr_addr_reg_bits_0 = _RAND_8[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  wr_data_1_valid = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  wr_data_1_bits = _RAND_10[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  wr_data_2_valid = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  wr_data_2_bits = _RAND_12[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  wr_addr_2 = _RAND_13[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  wr_data_final = _RAND_14[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  wr_addr_3 = _RAND_15[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  wr_valid_3 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_46 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_49 = _RAND_18[15:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(mem__T_43_en & mem__T_43_mask) begin
      mem[mem__T_43_addr] <= mem__T_43_data; // @[mem.scala 105:24]
    end
    mem_mem_output_en_pipe_0 <= rd_addr_reg_valid;
    if (rd_addr_reg_valid) begin
      mem_mem_output_addr_pipe_0 <= mem_rd_addr[2:0];
    end
    if (reset) begin
      rd_addr_reg_valid <= 1'h0;
    end else begin
      rd_addr_reg_valid <= io_rd_addr_valid;
    end
    if (reset) begin
      rd_addr_reg_bits_1 <= 16'h0;
    end else if (_T_14) begin
      rd_addr_reg_bits_1 <= 16'h0;
    end else if (_T_12) begin
      rd_addr_reg_bits_1 <= _T_11;
    end
    if (reset) begin
      rd_addr_reg_bits_0 <= 16'h0;
    end else if (_T_9) begin
      rd_addr_reg_bits_0 <= 16'h0;
    end else if (_T_7) begin
      rd_addr_reg_bits_0 <= _T_6;
    end
    if (reset) begin
      mem_req_valid <= 1'h0;
    end else begin
      mem_req_valid <= rd_addr_reg_valid;
    end
    if (reset) begin
      wr_addr_reg_bits_1 <= 16'h0;
    end else if (_T_30) begin
      wr_addr_reg_bits_1 <= 16'h0;
    end else if (_T_28) begin
      wr_addr_reg_bits_1 <= _T_27;
    end
    if (reset) begin
      wr_addr_reg_bits_0 <= 16'h0;
    end else if (_T_25) begin
      wr_addr_reg_bits_0 <= 16'h0;
    end else if (_T_23) begin
      wr_addr_reg_bits_0 <= _T_22;
    end
    if (reset) begin
      wr_data_1_valid <= 1'h0;
    end else begin
      wr_data_1_valid <= io_wr_data_valid;
    end
    if (reset) begin
      wr_data_1_bits <= 16'h0;
    end else begin
      wr_data_1_bits <= io_wr_data_bits;
    end
    if (reset) begin
      wr_data_2_valid <= 1'h0;
    end else begin
      wr_data_2_valid <= wr_data_1_valid;
    end
    if (reset) begin
      wr_data_2_bits <= 16'h0;
    end else begin
      wr_data_2_bits <= wr_data_1_bits;
    end
    if (reset) begin
      wr_addr_2 <= 16'h0;
    end else begin
      wr_addr_2 <= mem_wr_addr;
    end
    wr_data_final <= wr_data_2_bits;
    if (reset) begin
      wr_addr_3 <= 16'h0;
    end else begin
      wr_addr_3 <= wr_addr_2;
    end
    wr_valid_3 <= wr_data_2_valid;
    _T_46 <= mem_req_valid & mem_mem_output_data[16];
    if (mem_req_valid) begin
      _T_49 <= mem_mem_output_data[15:0];
    end else begin
      _T_49 <= 16'h0;
    end
  end
endmodule
module MemController(
  input         clock,
  input         reset,
  input         io_rd_valid,
  input         io_wr_valid,
  output        io_rd_data_valid,
  output [15:0] io_rd_data_bits,
  input         io_wr_data_valid,
  input  [15:0] io_wr_data_bits
);
  wire  MultiDimMem_clock; // @[mem.scala 32:19]
  wire  MultiDimMem_reset; // @[mem.scala 32:19]
  wire  MultiDimMem_io_rd_addr_valid; // @[mem.scala 32:19]
  wire [1:0] MultiDimMem_io_rd_addr_bits_0; // @[mem.scala 32:19]
  wire [1:0] MultiDimMem_io_rd_addr_bits_1; // @[mem.scala 32:19]
  wire  MultiDimMem_io_rd_data_valid; // @[mem.scala 32:19]
  wire [15:0] MultiDimMem_io_rd_data_bits; // @[mem.scala 32:19]
  wire [1:0] MultiDimMem_io_wr_addr_bits_0; // @[mem.scala 32:19]
  wire [1:0] MultiDimMem_io_wr_addr_bits_1; // @[mem.scala 32:19]
  wire  MultiDimMem_io_wr_data_valid; // @[mem.scala 32:19]
  wire [15:0] MultiDimMem_io_wr_data_bits; // @[mem.scala 32:19]
  wire  MultiDimTime_clock; // @[mem.scala 33:23]
  wire  MultiDimTime_reset; // @[mem.scala 33:23]
  wire  MultiDimTime_io_in; // @[mem.scala 33:23]
  wire [1:0] MultiDimTime_io_out_0; // @[mem.scala 33:23]
  wire [1:0] MultiDimTime_io_out_1; // @[mem.scala 33:23]
  wire [17:0] MultiDimTime_io_index_0; // @[mem.scala 33:23]
  wire [17:0] MultiDimTime_io_index_1; // @[mem.scala 33:23]
  wire  MultiDimTime_1_clock; // @[mem.scala 34:23]
  wire  MultiDimTime_1_reset; // @[mem.scala 34:23]
  wire  MultiDimTime_1_io_in; // @[mem.scala 34:23]
  wire [1:0] MultiDimTime_1_io_out_0; // @[mem.scala 34:23]
  wire [1:0] MultiDimTime_1_io_out_1; // @[mem.scala 34:23]
  wire [17:0] MultiDimTime_1_io_index_0; // @[mem.scala 34:23]
  wire [17:0] MultiDimTime_1_io_index_1; // @[mem.scala 34:23]
  MultiDimMem MultiDimMem ( // @[mem.scala 32:19]
    .clock(MultiDimMem_clock),
    .reset(MultiDimMem_reset),
    .io_rd_addr_valid(MultiDimMem_io_rd_addr_valid),
    .io_rd_addr_bits_0(MultiDimMem_io_rd_addr_bits_0),
    .io_rd_addr_bits_1(MultiDimMem_io_rd_addr_bits_1),
    .io_rd_data_valid(MultiDimMem_io_rd_data_valid),
    .io_rd_data_bits(MultiDimMem_io_rd_data_bits),
    .io_wr_addr_bits_0(MultiDimMem_io_wr_addr_bits_0),
    .io_wr_addr_bits_1(MultiDimMem_io_wr_addr_bits_1),
    .io_wr_data_valid(MultiDimMem_io_wr_data_valid),
    .io_wr_data_bits(MultiDimMem_io_wr_data_bits)
  );
  MultiDimTime MultiDimTime ( // @[mem.scala 33:23]
    .clock(MultiDimTime_clock),
    .reset(MultiDimTime_reset),
    .io_in(MultiDimTime_io_in),
    .io_out_0(MultiDimTime_io_out_0),
    .io_out_1(MultiDimTime_io_out_1),
    .io_index_0(MultiDimTime_io_index_0),
    .io_index_1(MultiDimTime_io_index_1)
  );
  MultiDimTime MultiDimTime_1 ( // @[mem.scala 34:23]
    .clock(MultiDimTime_1_clock),
    .reset(MultiDimTime_1_reset),
    .io_in(MultiDimTime_1_io_in),
    .io_out_0(MultiDimTime_1_io_out_0),
    .io_out_1(MultiDimTime_1_io_out_1),
    .io_index_0(MultiDimTime_1_io_index_0),
    .io_index_1(MultiDimTime_1_io_index_1)
  );
  assign io_rd_data_valid = MultiDimMem_io_rd_data_valid; // @[mem.scala 52:14]
  assign io_rd_data_bits = MultiDimMem_io_rd_data_bits; // @[mem.scala 52:14]
  assign MultiDimMem_clock = clock;
  assign MultiDimMem_reset = reset;
  assign MultiDimMem_io_rd_addr_valid = io_rd_valid; // @[mem.scala 49:21]
  assign MultiDimMem_io_rd_addr_bits_0 = MultiDimTime_1_io_out_0; // @[mem.scala 48:20]
  assign MultiDimMem_io_rd_addr_bits_1 = MultiDimTime_1_io_out_1; // @[mem.scala 48:20]
  assign MultiDimMem_io_wr_addr_bits_0 = MultiDimTime_io_out_0; // @[mem.scala 44:20]
  assign MultiDimMem_io_wr_addr_bits_1 = MultiDimTime_io_out_1; // @[mem.scala 44:20]
  assign MultiDimMem_io_wr_data_valid = io_wr_data_valid; // @[mem.scala 53:15]
  assign MultiDimMem_io_wr_data_bits = io_wr_data_bits; // @[mem.scala 53:15]
  assign MultiDimTime_clock = clock;
  assign MultiDimTime_reset = reset;
  assign MultiDimTime_io_in = io_wr_valid; // @[mem.scala 43:14]
  assign MultiDimTime_1_clock = clock;
  assign MultiDimTime_1_reset = reset;
  assign MultiDimTime_1_io_in = io_rd_valid; // @[mem.scala 47:14]
endmodule
module PEArray(
  input         clock,
  input         reset,
  input         io_data_2_in_0_valid,
  input         io_data_2_in_0_bits_valid,
  input  [15:0] io_data_2_in_0_bits_bits,
  input         io_data_2_in_1_valid,
  input         io_data_2_in_1_bits_valid,
  input  [15:0] io_data_2_in_1_bits_bits,
  input         io_data_2_in_2_valid,
  input         io_data_2_in_2_bits_valid,
  input  [15:0] io_data_2_in_2_bits_bits,
  input         io_data_2_in_3_valid,
  input         io_data_2_in_3_bits_valid,
  input  [15:0] io_data_2_in_3_bits_bits,
  input         io_data_2_in_4_valid,
  input         io_data_2_in_4_bits_valid,
  input  [15:0] io_data_2_in_4_bits_bits,
  input         io_data_2_in_5_valid,
  input         io_data_2_in_5_bits_valid,
  input  [15:0] io_data_2_in_5_bits_bits,
  input         io_data_2_in_6_valid,
  input         io_data_2_in_6_bits_valid,
  input  [15:0] io_data_2_in_6_bits_bits,
  input         io_data_2_in_7_valid,
  input         io_data_2_in_7_bits_valid,
  input  [15:0] io_data_2_in_7_bits_bits,
  input         io_data_1_in_0_valid,
  input         io_data_1_in_0_bits_valid,
  input  [15:0] io_data_1_in_0_bits_bits,
  input         io_data_1_in_1_valid,
  input         io_data_1_in_1_bits_valid,
  input  [15:0] io_data_1_in_1_bits_bits,
  input         io_data_1_in_2_valid,
  input         io_data_1_in_2_bits_valid,
  input  [15:0] io_data_1_in_2_bits_bits,
  input         io_data_1_in_3_valid,
  input         io_data_1_in_3_bits_valid,
  input  [15:0] io_data_1_in_3_bits_bits,
  input         io_data_1_in_4_valid,
  input         io_data_1_in_4_bits_valid,
  input  [15:0] io_data_1_in_4_bits_bits,
  input         io_data_1_in_5_valid,
  input         io_data_1_in_5_bits_valid,
  input  [15:0] io_data_1_in_5_bits_bits,
  input         io_data_1_in_6_valid,
  input         io_data_1_in_6_bits_valid,
  input  [15:0] io_data_1_in_6_bits_bits,
  input         io_data_1_in_7_valid,
  input         io_data_1_in_7_bits_valid,
  input  [15:0] io_data_1_in_7_bits_bits,
  output        io_data_0_out_0_valid,
  output [15:0] io_data_0_out_0_bits,
  output        io_data_0_out_1_valid,
  output [15:0] io_data_0_out_1_bits,
  output        io_data_0_out_2_valid,
  output [15:0] io_data_0_out_2_bits,
  output        io_data_0_out_3_valid,
  output [15:0] io_data_0_out_3_bits,
  output        io_data_0_out_4_valid,
  output [15:0] io_data_0_out_4_bits,
  output        io_data_0_out_5_valid,
  output [15:0] io_data_0_out_5_bits,
  output        io_data_0_out_6_valid,
  output [15:0] io_data_0_out_6_bits,
  output        io_data_0_out_7_valid,
  output [15:0] io_data_0_out_7_bits,
  input         io_exec_valid,
  input         io_out_valid
);
  wire  MultiDimTime_clock; // @[pearray.scala 63:25]
  wire  MultiDimTime_reset; // @[pearray.scala 63:25]
  wire  MultiDimTime_io_in; // @[pearray.scala 63:25]
  wire [1:0] MultiDimTime_io_out_0; // @[pearray.scala 63:25]
  wire [1:0] MultiDimTime_io_out_1; // @[pearray.scala 63:25]
  wire [17:0] MultiDimTime_io_index_0; // @[pearray.scala 63:25]
  wire [17:0] MultiDimTime_io_index_1; // @[pearray.scala 63:25]
  wire  PE_clock; // @[pearray.scala 103:13]
  wire  PE_reset; // @[pearray.scala 103:13]
  wire  PE_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_1_clock; // @[pearray.scala 103:13]
  wire  PE_1_reset; // @[pearray.scala 103:13]
  wire  PE_1_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_1_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_1_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_1_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_1_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_1_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_1_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_1_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_1_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_1_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_1_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_1_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_1_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_2_clock; // @[pearray.scala 103:13]
  wire  PE_2_reset; // @[pearray.scala 103:13]
  wire  PE_2_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_2_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_2_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_2_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_2_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_2_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_2_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_2_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_2_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_2_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_2_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_2_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_2_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_3_clock; // @[pearray.scala 103:13]
  wire  PE_3_reset; // @[pearray.scala 103:13]
  wire  PE_3_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_3_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_3_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_3_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_3_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_3_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_3_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_3_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_3_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_3_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_3_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_3_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_3_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_4_clock; // @[pearray.scala 103:13]
  wire  PE_4_reset; // @[pearray.scala 103:13]
  wire  PE_4_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_4_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_4_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_4_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_4_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_4_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_4_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_4_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_4_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_4_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_4_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_4_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_4_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_5_clock; // @[pearray.scala 103:13]
  wire  PE_5_reset; // @[pearray.scala 103:13]
  wire  PE_5_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_5_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_5_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_5_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_5_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_5_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_5_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_5_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_5_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_5_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_5_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_5_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_5_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_6_clock; // @[pearray.scala 103:13]
  wire  PE_6_reset; // @[pearray.scala 103:13]
  wire  PE_6_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_6_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_6_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_6_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_6_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_6_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_6_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_6_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_6_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_6_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_6_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_6_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_6_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_7_clock; // @[pearray.scala 103:13]
  wire  PE_7_reset; // @[pearray.scala 103:13]
  wire  PE_7_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_7_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_7_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_7_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_7_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_7_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_7_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_7_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_7_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_7_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_7_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_7_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_7_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_8_clock; // @[pearray.scala 103:13]
  wire  PE_8_reset; // @[pearray.scala 103:13]
  wire  PE_8_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_8_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_8_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_8_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_8_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_8_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_8_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_8_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_8_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_8_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_8_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_8_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_8_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_9_clock; // @[pearray.scala 103:13]
  wire  PE_9_reset; // @[pearray.scala 103:13]
  wire  PE_9_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_9_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_9_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_9_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_9_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_9_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_9_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_9_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_9_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_9_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_9_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_9_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_9_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_10_clock; // @[pearray.scala 103:13]
  wire  PE_10_reset; // @[pearray.scala 103:13]
  wire  PE_10_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_10_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_10_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_10_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_10_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_10_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_10_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_10_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_10_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_10_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_10_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_10_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_10_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_11_clock; // @[pearray.scala 103:13]
  wire  PE_11_reset; // @[pearray.scala 103:13]
  wire  PE_11_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_11_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_11_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_11_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_11_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_11_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_11_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_11_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_11_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_11_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_11_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_11_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_11_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_12_clock; // @[pearray.scala 103:13]
  wire  PE_12_reset; // @[pearray.scala 103:13]
  wire  PE_12_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_12_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_12_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_12_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_12_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_12_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_12_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_12_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_12_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_12_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_12_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_12_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_12_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_13_clock; // @[pearray.scala 103:13]
  wire  PE_13_reset; // @[pearray.scala 103:13]
  wire  PE_13_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_13_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_13_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_13_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_13_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_13_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_13_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_13_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_13_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_13_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_13_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_13_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_13_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_14_clock; // @[pearray.scala 103:13]
  wire  PE_14_reset; // @[pearray.scala 103:13]
  wire  PE_14_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_14_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_14_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_14_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_14_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_14_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_14_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_14_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_14_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_14_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_14_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_14_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_14_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_15_clock; // @[pearray.scala 103:13]
  wire  PE_15_reset; // @[pearray.scala 103:13]
  wire  PE_15_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_15_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_15_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_15_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_15_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_15_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_15_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_15_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_15_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_15_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_15_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_15_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_15_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_16_clock; // @[pearray.scala 103:13]
  wire  PE_16_reset; // @[pearray.scala 103:13]
  wire  PE_16_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_16_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_16_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_16_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_16_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_16_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_16_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_16_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_16_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_16_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_16_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_16_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_16_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_17_clock; // @[pearray.scala 103:13]
  wire  PE_17_reset; // @[pearray.scala 103:13]
  wire  PE_17_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_17_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_17_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_17_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_17_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_17_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_17_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_17_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_17_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_17_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_17_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_17_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_17_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_18_clock; // @[pearray.scala 103:13]
  wire  PE_18_reset; // @[pearray.scala 103:13]
  wire  PE_18_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_18_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_18_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_18_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_18_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_18_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_18_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_18_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_18_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_18_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_18_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_18_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_18_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_19_clock; // @[pearray.scala 103:13]
  wire  PE_19_reset; // @[pearray.scala 103:13]
  wire  PE_19_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_19_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_19_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_19_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_19_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_19_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_19_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_19_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_19_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_19_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_19_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_19_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_19_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_20_clock; // @[pearray.scala 103:13]
  wire  PE_20_reset; // @[pearray.scala 103:13]
  wire  PE_20_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_20_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_20_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_20_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_20_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_20_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_20_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_20_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_20_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_20_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_20_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_20_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_20_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_21_clock; // @[pearray.scala 103:13]
  wire  PE_21_reset; // @[pearray.scala 103:13]
  wire  PE_21_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_21_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_21_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_21_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_21_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_21_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_21_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_21_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_21_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_21_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_21_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_21_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_21_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_22_clock; // @[pearray.scala 103:13]
  wire  PE_22_reset; // @[pearray.scala 103:13]
  wire  PE_22_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_22_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_22_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_22_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_22_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_22_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_22_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_22_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_22_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_22_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_22_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_22_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_22_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_23_clock; // @[pearray.scala 103:13]
  wire  PE_23_reset; // @[pearray.scala 103:13]
  wire  PE_23_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_23_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_23_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_23_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_23_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_23_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_23_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_23_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_23_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_23_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_23_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_23_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_23_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_24_clock; // @[pearray.scala 103:13]
  wire  PE_24_reset; // @[pearray.scala 103:13]
  wire  PE_24_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_24_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_24_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_24_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_24_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_24_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_24_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_24_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_24_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_24_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_24_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_24_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_24_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_25_clock; // @[pearray.scala 103:13]
  wire  PE_25_reset; // @[pearray.scala 103:13]
  wire  PE_25_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_25_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_25_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_25_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_25_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_25_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_25_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_25_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_25_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_25_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_25_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_25_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_25_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_26_clock; // @[pearray.scala 103:13]
  wire  PE_26_reset; // @[pearray.scala 103:13]
  wire  PE_26_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_26_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_26_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_26_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_26_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_26_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_26_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_26_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_26_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_26_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_26_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_26_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_26_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_27_clock; // @[pearray.scala 103:13]
  wire  PE_27_reset; // @[pearray.scala 103:13]
  wire  PE_27_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_27_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_27_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_27_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_27_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_27_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_27_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_27_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_27_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_27_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_27_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_27_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_27_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_28_clock; // @[pearray.scala 103:13]
  wire  PE_28_reset; // @[pearray.scala 103:13]
  wire  PE_28_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_28_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_28_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_28_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_28_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_28_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_28_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_28_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_28_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_28_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_28_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_28_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_28_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_29_clock; // @[pearray.scala 103:13]
  wire  PE_29_reset; // @[pearray.scala 103:13]
  wire  PE_29_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_29_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_29_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_29_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_29_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_29_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_29_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_29_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_29_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_29_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_29_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_29_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_29_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_30_clock; // @[pearray.scala 103:13]
  wire  PE_30_reset; // @[pearray.scala 103:13]
  wire  PE_30_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_30_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_30_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_30_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_30_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_30_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_30_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_30_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_30_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_30_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_30_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_30_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_30_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_31_clock; // @[pearray.scala 103:13]
  wire  PE_31_reset; // @[pearray.scala 103:13]
  wire  PE_31_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_31_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_31_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_31_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_31_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_31_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_31_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_31_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_31_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_31_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_31_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_31_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_31_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_32_clock; // @[pearray.scala 103:13]
  wire  PE_32_reset; // @[pearray.scala 103:13]
  wire  PE_32_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_32_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_32_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_32_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_32_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_32_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_32_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_32_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_32_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_32_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_32_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_32_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_32_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_33_clock; // @[pearray.scala 103:13]
  wire  PE_33_reset; // @[pearray.scala 103:13]
  wire  PE_33_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_33_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_33_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_33_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_33_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_33_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_33_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_33_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_33_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_33_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_33_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_33_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_33_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_34_clock; // @[pearray.scala 103:13]
  wire  PE_34_reset; // @[pearray.scala 103:13]
  wire  PE_34_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_34_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_34_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_34_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_34_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_34_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_34_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_34_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_34_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_34_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_34_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_34_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_34_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_35_clock; // @[pearray.scala 103:13]
  wire  PE_35_reset; // @[pearray.scala 103:13]
  wire  PE_35_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_35_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_35_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_35_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_35_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_35_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_35_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_35_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_35_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_35_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_35_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_35_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_35_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_36_clock; // @[pearray.scala 103:13]
  wire  PE_36_reset; // @[pearray.scala 103:13]
  wire  PE_36_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_36_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_36_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_36_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_36_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_36_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_36_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_36_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_36_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_36_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_36_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_36_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_36_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_37_clock; // @[pearray.scala 103:13]
  wire  PE_37_reset; // @[pearray.scala 103:13]
  wire  PE_37_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_37_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_37_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_37_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_37_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_37_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_37_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_37_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_37_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_37_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_37_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_37_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_37_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_38_clock; // @[pearray.scala 103:13]
  wire  PE_38_reset; // @[pearray.scala 103:13]
  wire  PE_38_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_38_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_38_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_38_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_38_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_38_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_38_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_38_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_38_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_38_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_38_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_38_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_38_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_39_clock; // @[pearray.scala 103:13]
  wire  PE_39_reset; // @[pearray.scala 103:13]
  wire  PE_39_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_39_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_39_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_39_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_39_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_39_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_39_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_39_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_39_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_39_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_39_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_39_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_39_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_40_clock; // @[pearray.scala 103:13]
  wire  PE_40_reset; // @[pearray.scala 103:13]
  wire  PE_40_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_40_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_40_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_40_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_40_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_40_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_40_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_40_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_40_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_40_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_40_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_40_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_40_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_41_clock; // @[pearray.scala 103:13]
  wire  PE_41_reset; // @[pearray.scala 103:13]
  wire  PE_41_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_41_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_41_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_41_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_41_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_41_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_41_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_41_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_41_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_41_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_41_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_41_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_41_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_42_clock; // @[pearray.scala 103:13]
  wire  PE_42_reset; // @[pearray.scala 103:13]
  wire  PE_42_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_42_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_42_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_42_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_42_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_42_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_42_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_42_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_42_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_42_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_42_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_42_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_42_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_43_clock; // @[pearray.scala 103:13]
  wire  PE_43_reset; // @[pearray.scala 103:13]
  wire  PE_43_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_43_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_43_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_43_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_43_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_43_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_43_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_43_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_43_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_43_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_43_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_43_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_43_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_44_clock; // @[pearray.scala 103:13]
  wire  PE_44_reset; // @[pearray.scala 103:13]
  wire  PE_44_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_44_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_44_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_44_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_44_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_44_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_44_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_44_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_44_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_44_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_44_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_44_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_44_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_45_clock; // @[pearray.scala 103:13]
  wire  PE_45_reset; // @[pearray.scala 103:13]
  wire  PE_45_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_45_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_45_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_45_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_45_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_45_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_45_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_45_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_45_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_45_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_45_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_45_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_45_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_46_clock; // @[pearray.scala 103:13]
  wire  PE_46_reset; // @[pearray.scala 103:13]
  wire  PE_46_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_46_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_46_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_46_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_46_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_46_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_46_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_46_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_46_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_46_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_46_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_46_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_46_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_47_clock; // @[pearray.scala 103:13]
  wire  PE_47_reset; // @[pearray.scala 103:13]
  wire  PE_47_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_47_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_47_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_47_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_47_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_47_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_47_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_47_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_47_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_47_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_47_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_47_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_47_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_48_clock; // @[pearray.scala 103:13]
  wire  PE_48_reset; // @[pearray.scala 103:13]
  wire  PE_48_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_48_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_48_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_48_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_48_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_48_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_48_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_48_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_48_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_48_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_48_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_48_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_48_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_49_clock; // @[pearray.scala 103:13]
  wire  PE_49_reset; // @[pearray.scala 103:13]
  wire  PE_49_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_49_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_49_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_49_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_49_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_49_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_49_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_49_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_49_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_49_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_49_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_49_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_49_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_50_clock; // @[pearray.scala 103:13]
  wire  PE_50_reset; // @[pearray.scala 103:13]
  wire  PE_50_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_50_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_50_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_50_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_50_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_50_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_50_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_50_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_50_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_50_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_50_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_50_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_50_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_51_clock; // @[pearray.scala 103:13]
  wire  PE_51_reset; // @[pearray.scala 103:13]
  wire  PE_51_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_51_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_51_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_51_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_51_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_51_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_51_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_51_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_51_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_51_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_51_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_51_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_51_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_52_clock; // @[pearray.scala 103:13]
  wire  PE_52_reset; // @[pearray.scala 103:13]
  wire  PE_52_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_52_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_52_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_52_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_52_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_52_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_52_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_52_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_52_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_52_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_52_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_52_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_52_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_53_clock; // @[pearray.scala 103:13]
  wire  PE_53_reset; // @[pearray.scala 103:13]
  wire  PE_53_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_53_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_53_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_53_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_53_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_53_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_53_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_53_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_53_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_53_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_53_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_53_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_53_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_54_clock; // @[pearray.scala 103:13]
  wire  PE_54_reset; // @[pearray.scala 103:13]
  wire  PE_54_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_54_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_54_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_54_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_54_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_54_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_54_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_54_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_54_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_54_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_54_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_54_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_54_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_55_clock; // @[pearray.scala 103:13]
  wire  PE_55_reset; // @[pearray.scala 103:13]
  wire  PE_55_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_55_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_55_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_55_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_55_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_55_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_55_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_55_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_55_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_55_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_55_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_55_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_55_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_56_clock; // @[pearray.scala 103:13]
  wire  PE_56_reset; // @[pearray.scala 103:13]
  wire  PE_56_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_56_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_56_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_56_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_56_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_56_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_56_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_56_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_56_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_56_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_56_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_56_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_56_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_57_clock; // @[pearray.scala 103:13]
  wire  PE_57_reset; // @[pearray.scala 103:13]
  wire  PE_57_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_57_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_57_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_57_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_57_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_57_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_57_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_57_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_57_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_57_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_57_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_57_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_57_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_58_clock; // @[pearray.scala 103:13]
  wire  PE_58_reset; // @[pearray.scala 103:13]
  wire  PE_58_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_58_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_58_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_58_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_58_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_58_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_58_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_58_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_58_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_58_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_58_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_58_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_58_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_59_clock; // @[pearray.scala 103:13]
  wire  PE_59_reset; // @[pearray.scala 103:13]
  wire  PE_59_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_59_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_59_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_59_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_59_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_59_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_59_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_59_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_59_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_59_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_59_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_59_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_59_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_60_clock; // @[pearray.scala 103:13]
  wire  PE_60_reset; // @[pearray.scala 103:13]
  wire  PE_60_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_60_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_60_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_60_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_60_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_60_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_60_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_60_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_60_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_60_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_60_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_60_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_60_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_61_clock; // @[pearray.scala 103:13]
  wire  PE_61_reset; // @[pearray.scala 103:13]
  wire  PE_61_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_61_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_61_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_61_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_61_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_61_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_61_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_61_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_61_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_61_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_61_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_61_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_61_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_62_clock; // @[pearray.scala 103:13]
  wire  PE_62_reset; // @[pearray.scala 103:13]
  wire  PE_62_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_62_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_62_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_62_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_62_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_62_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_62_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_62_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_62_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_62_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_62_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_62_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_62_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PE_63_clock; // @[pearray.scala 103:13]
  wire  PE_63_reset; // @[pearray.scala 103:13]
  wire  PE_63_io_data_2_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_63_io_data_2_in_bits; // @[pearray.scala 103:13]
  wire  PE_63_io_data_2_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_63_io_data_2_out_bits; // @[pearray.scala 103:13]
  wire  PE_63_io_data_1_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_63_io_data_1_in_bits; // @[pearray.scala 103:13]
  wire  PE_63_io_data_1_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_63_io_data_1_out_bits; // @[pearray.scala 103:13]
  wire  PE_63_io_data_0_in_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_63_io_data_0_in_bits; // @[pearray.scala 103:13]
  wire  PE_63_io_data_0_out_valid; // @[pearray.scala 103:13]
  wire [15:0] PE_63_io_data_0_out_bits; // @[pearray.scala 103:13]
  wire  PE_63_io_sig_stat2trans; // @[pearray.scala 103:13]
  wire  PENetwork_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_io_to_pes_7_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_io_to_pes_7_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_1_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_1_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_1_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_1_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_1_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_1_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_1_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_1_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_1_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_1_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_1_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_1_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_1_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_1_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_1_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_1_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_1_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_1_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_1_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_1_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_1_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_1_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_1_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_1_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_1_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_1_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_1_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_1_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_1_io_to_pes_7_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_1_io_to_pes_7_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_1_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_1_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_2_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_2_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_2_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_2_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_2_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_2_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_2_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_2_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_2_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_2_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_2_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_2_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_2_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_2_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_2_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_2_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_2_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_2_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_2_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_2_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_2_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_2_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_2_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_2_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_2_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_2_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_2_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_2_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_2_io_to_pes_7_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_2_io_to_pes_7_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_2_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_2_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_3_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_3_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_3_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_3_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_3_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_3_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_3_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_3_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_3_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_3_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_3_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_3_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_3_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_3_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_3_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_3_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_3_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_3_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_3_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_3_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_3_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_3_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_3_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_3_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_3_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_3_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_3_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_3_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_3_io_to_pes_7_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_3_io_to_pes_7_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_3_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_3_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_4_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_4_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_4_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_4_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_4_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_4_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_4_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_4_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_4_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_4_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_4_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_4_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_4_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_4_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_4_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_4_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_4_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_4_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_4_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_4_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_4_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_4_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_4_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_4_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_4_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_4_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_4_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_4_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_4_io_to_pes_7_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_4_io_to_pes_7_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_4_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_4_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_5_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_5_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_5_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_5_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_5_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_5_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_5_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_5_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_5_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_5_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_5_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_5_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_5_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_5_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_5_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_5_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_5_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_5_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_5_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_5_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_5_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_5_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_5_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_5_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_5_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_5_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_5_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_5_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_5_io_to_pes_7_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_5_io_to_pes_7_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_5_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_5_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_6_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_6_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_6_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_6_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_6_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_6_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_6_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_6_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_6_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_6_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_6_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_6_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_6_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_6_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_6_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_6_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_6_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_6_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_6_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_6_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_6_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_6_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_6_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_6_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_6_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_6_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_6_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_6_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_6_io_to_pes_7_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_6_io_to_pes_7_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_6_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_6_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_7_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_7_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_7_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_7_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_7_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_7_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_7_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_7_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_7_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_7_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_7_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_7_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_7_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_7_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_7_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_7_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_7_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_7_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_7_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_7_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_7_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_7_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_7_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_7_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_7_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_7_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_7_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_7_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_7_io_to_pes_7_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_7_io_to_pes_7_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_7_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_7_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_8_io_to_pes_0_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_8_io_to_pes_0_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_8_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_8_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_8_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_8_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_8_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_8_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_8_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_8_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_8_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_8_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_8_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_8_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_8_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_8_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_8_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_8_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_8_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_8_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_8_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_8_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_8_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_8_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_8_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_8_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_8_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_8_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_8_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_8_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_8_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_8_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_9_io_to_pes_0_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_9_io_to_pes_0_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_9_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_9_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_9_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_9_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_9_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_9_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_9_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_9_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_9_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_9_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_9_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_9_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_9_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_9_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_9_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_9_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_9_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_9_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_9_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_9_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_9_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_9_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_9_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_9_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_9_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_9_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_9_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_9_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_9_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_9_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_10_io_to_pes_0_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_10_io_to_pes_0_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_10_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_10_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_10_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_10_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_10_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_10_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_10_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_10_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_10_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_10_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_10_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_10_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_10_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_10_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_10_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_10_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_10_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_10_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_10_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_10_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_10_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_10_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_10_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_10_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_10_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_10_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_10_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_10_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_10_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_10_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_11_io_to_pes_0_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_11_io_to_pes_0_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_11_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_11_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_11_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_11_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_11_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_11_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_11_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_11_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_11_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_11_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_11_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_11_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_11_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_11_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_11_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_11_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_11_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_11_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_11_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_11_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_11_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_11_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_11_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_11_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_11_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_11_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_11_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_11_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_11_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_11_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_12_io_to_pes_0_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_12_io_to_pes_0_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_12_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_12_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_12_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_12_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_12_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_12_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_12_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_12_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_12_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_12_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_12_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_12_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_12_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_12_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_12_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_12_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_12_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_12_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_12_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_12_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_12_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_12_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_12_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_12_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_12_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_12_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_12_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_12_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_12_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_12_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_13_io_to_pes_0_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_13_io_to_pes_0_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_13_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_13_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_13_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_13_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_13_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_13_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_13_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_13_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_13_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_13_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_13_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_13_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_13_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_13_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_13_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_13_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_13_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_13_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_13_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_13_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_13_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_13_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_13_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_13_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_13_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_13_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_13_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_13_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_13_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_13_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_14_io_to_pes_0_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_14_io_to_pes_0_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_14_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_14_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_14_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_14_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_14_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_14_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_14_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_14_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_14_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_14_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_14_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_14_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_14_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_14_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_14_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_14_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_14_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_14_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_14_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_14_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_14_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_14_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_14_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_14_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_14_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_14_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_14_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_14_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_14_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_14_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_15_io_to_pes_0_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_15_io_to_pes_0_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_15_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_15_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_15_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_15_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_15_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_15_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_15_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_15_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_15_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_15_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_15_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_15_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_15_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_15_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_15_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_15_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_15_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_15_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_15_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_15_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_15_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_15_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_15_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_15_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_15_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_15_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_15_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_15_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_15_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_15_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_16_io_to_pes_0_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_16_io_to_pes_0_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_16_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_16_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_16_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_16_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_16_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_16_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_16_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_16_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_16_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_16_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_16_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_16_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_16_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_16_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_16_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_16_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_16_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_16_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_16_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_16_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_16_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_16_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_16_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_16_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_16_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_16_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_16_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_16_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_16_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_16_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_17_io_to_pes_0_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_17_io_to_pes_0_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_17_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_17_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_17_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_17_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_17_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_17_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_17_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_17_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_17_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_17_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_17_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_17_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_17_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_17_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_17_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_17_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_17_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_17_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_17_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_17_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_17_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_17_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_17_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_17_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_17_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_17_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_17_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_17_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_17_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_17_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_18_io_to_pes_0_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_18_io_to_pes_0_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_18_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_18_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_18_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_18_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_18_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_18_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_18_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_18_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_18_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_18_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_18_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_18_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_18_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_18_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_18_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_18_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_18_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_18_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_18_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_18_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_18_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_18_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_18_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_18_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_18_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_18_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_18_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_18_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_18_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_18_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_19_io_to_pes_0_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_19_io_to_pes_0_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_19_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_19_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_19_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_19_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_19_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_19_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_19_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_19_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_19_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_19_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_19_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_19_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_19_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_19_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_19_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_19_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_19_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_19_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_19_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_19_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_19_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_19_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_19_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_19_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_19_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_19_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_19_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_19_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_19_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_19_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_20_io_to_pes_0_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_20_io_to_pes_0_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_20_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_20_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_20_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_20_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_20_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_20_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_20_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_20_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_20_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_20_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_20_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_20_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_20_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_20_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_20_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_20_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_20_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_20_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_20_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_20_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_20_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_20_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_20_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_20_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_20_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_20_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_20_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_20_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_20_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_20_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_21_io_to_pes_0_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_21_io_to_pes_0_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_21_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_21_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_21_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_21_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_21_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_21_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_21_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_21_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_21_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_21_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_21_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_21_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_21_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_21_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_21_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_21_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_21_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_21_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_21_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_21_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_21_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_21_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_21_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_21_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_21_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_21_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_21_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_21_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_21_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_21_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_22_io_to_pes_0_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_22_io_to_pes_0_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_22_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_22_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_22_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_22_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_22_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_22_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_22_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_22_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_22_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_22_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_22_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_22_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_22_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_22_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_22_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_22_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_22_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_22_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_22_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_22_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_22_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_22_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_22_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_22_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_22_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_22_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_22_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_22_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_22_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_22_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  PENetwork_23_io_to_pes_0_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_23_io_to_pes_0_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_23_io_to_pes_0_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_23_io_to_pes_0_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_23_io_to_pes_1_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_23_io_to_pes_1_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_23_io_to_pes_1_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_23_io_to_pes_1_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_23_io_to_pes_2_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_23_io_to_pes_2_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_23_io_to_pes_2_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_23_io_to_pes_2_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_23_io_to_pes_3_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_23_io_to_pes_3_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_23_io_to_pes_3_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_23_io_to_pes_3_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_23_io_to_pes_4_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_23_io_to_pes_4_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_23_io_to_pes_4_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_23_io_to_pes_4_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_23_io_to_pes_5_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_23_io_to_pes_5_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_23_io_to_pes_5_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_23_io_to_pes_5_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_23_io_to_pes_6_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_23_io_to_pes_6_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_23_io_to_pes_6_out_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_23_io_to_pes_6_out_bits; // @[pearray.scala 137:13]
  wire  PENetwork_23_io_to_pes_7_in_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_23_io_to_pes_7_in_bits; // @[pearray.scala 137:13]
  wire  PENetwork_23_io_to_mem_valid; // @[pearray.scala 137:13]
  wire [15:0] PENetwork_23_io_to_mem_bits; // @[pearray.scala 137:13]
  wire  MemController_clock; // @[pearray.scala 211:15]
  wire  MemController_reset; // @[pearray.scala 211:15]
  wire  MemController_io_rd_valid; // @[pearray.scala 211:15]
  wire  MemController_io_wr_valid; // @[pearray.scala 211:15]
  wire  MemController_io_rd_data_valid; // @[pearray.scala 211:15]
  wire [15:0] MemController_io_rd_data_bits; // @[pearray.scala 211:15]
  wire  MemController_io_wr_data_valid; // @[pearray.scala 211:15]
  wire [15:0] MemController_io_wr_data_bits; // @[pearray.scala 211:15]
  wire  MemController_1_clock; // @[pearray.scala 211:15]
  wire  MemController_1_reset; // @[pearray.scala 211:15]
  wire  MemController_1_io_rd_valid; // @[pearray.scala 211:15]
  wire  MemController_1_io_wr_valid; // @[pearray.scala 211:15]
  wire  MemController_1_io_rd_data_valid; // @[pearray.scala 211:15]
  wire [15:0] MemController_1_io_rd_data_bits; // @[pearray.scala 211:15]
  wire  MemController_1_io_wr_data_valid; // @[pearray.scala 211:15]
  wire [15:0] MemController_1_io_wr_data_bits; // @[pearray.scala 211:15]
  wire  MemController_2_clock; // @[pearray.scala 211:15]
  wire  MemController_2_reset; // @[pearray.scala 211:15]
  wire  MemController_2_io_rd_valid; // @[pearray.scala 211:15]
  wire  MemController_2_io_wr_valid; // @[pearray.scala 211:15]
  wire  MemController_2_io_rd_data_valid; // @[pearray.scala 211:15]
  wire [15:0] MemController_2_io_rd_data_bits; // @[pearray.scala 211:15]
  wire  MemController_2_io_wr_data_valid; // @[pearray.scala 211:15]
  wire [15:0] MemController_2_io_wr_data_bits; // @[pearray.scala 211:15]
  wire  MemController_3_clock; // @[pearray.scala 211:15]
  wire  MemController_3_reset; // @[pearray.scala 211:15]
  wire  MemController_3_io_rd_valid; // @[pearray.scala 211:15]
  wire  MemController_3_io_wr_valid; // @[pearray.scala 211:15]
  wire  MemController_3_io_rd_data_valid; // @[pearray.scala 211:15]
  wire [15:0] MemController_3_io_rd_data_bits; // @[pearray.scala 211:15]
  wire  MemController_3_io_wr_data_valid; // @[pearray.scala 211:15]
  wire [15:0] MemController_3_io_wr_data_bits; // @[pearray.scala 211:15]
  wire  MemController_4_clock; // @[pearray.scala 211:15]
  wire  MemController_4_reset; // @[pearray.scala 211:15]
  wire  MemController_4_io_rd_valid; // @[pearray.scala 211:15]
  wire  MemController_4_io_wr_valid; // @[pearray.scala 211:15]
  wire  MemController_4_io_rd_data_valid; // @[pearray.scala 211:15]
  wire [15:0] MemController_4_io_rd_data_bits; // @[pearray.scala 211:15]
  wire  MemController_4_io_wr_data_valid; // @[pearray.scala 211:15]
  wire [15:0] MemController_4_io_wr_data_bits; // @[pearray.scala 211:15]
  wire  MemController_5_clock; // @[pearray.scala 211:15]
  wire  MemController_5_reset; // @[pearray.scala 211:15]
  wire  MemController_5_io_rd_valid; // @[pearray.scala 211:15]
  wire  MemController_5_io_wr_valid; // @[pearray.scala 211:15]
  wire  MemController_5_io_rd_data_valid; // @[pearray.scala 211:15]
  wire [15:0] MemController_5_io_rd_data_bits; // @[pearray.scala 211:15]
  wire  MemController_5_io_wr_data_valid; // @[pearray.scala 211:15]
  wire [15:0] MemController_5_io_wr_data_bits; // @[pearray.scala 211:15]
  wire  MemController_6_clock; // @[pearray.scala 211:15]
  wire  MemController_6_reset; // @[pearray.scala 211:15]
  wire  MemController_6_io_rd_valid; // @[pearray.scala 211:15]
  wire  MemController_6_io_wr_valid; // @[pearray.scala 211:15]
  wire  MemController_6_io_rd_data_valid; // @[pearray.scala 211:15]
  wire [15:0] MemController_6_io_rd_data_bits; // @[pearray.scala 211:15]
  wire  MemController_6_io_wr_data_valid; // @[pearray.scala 211:15]
  wire [15:0] MemController_6_io_wr_data_bits; // @[pearray.scala 211:15]
  wire  MemController_7_clock; // @[pearray.scala 211:15]
  wire  MemController_7_reset; // @[pearray.scala 211:15]
  wire  MemController_7_io_rd_valid; // @[pearray.scala 211:15]
  wire  MemController_7_io_wr_valid; // @[pearray.scala 211:15]
  wire  MemController_7_io_rd_data_valid; // @[pearray.scala 211:15]
  wire [15:0] MemController_7_io_rd_data_bits; // @[pearray.scala 211:15]
  wire  MemController_7_io_wr_data_valid; // @[pearray.scala 211:15]
  wire [15:0] MemController_7_io_wr_data_bits; // @[pearray.scala 211:15]
  wire  MemController_8_clock; // @[pearray.scala 209:15]
  wire  MemController_8_reset; // @[pearray.scala 209:15]
  wire  MemController_8_io_rd_valid; // @[pearray.scala 209:15]
  wire  MemController_8_io_wr_valid; // @[pearray.scala 209:15]
  wire  MemController_8_io_rd_data_valid; // @[pearray.scala 209:15]
  wire [15:0] MemController_8_io_rd_data_bits; // @[pearray.scala 209:15]
  wire  MemController_8_io_wr_data_valid; // @[pearray.scala 209:15]
  wire [15:0] MemController_8_io_wr_data_bits; // @[pearray.scala 209:15]
  wire  MemController_9_clock; // @[pearray.scala 209:15]
  wire  MemController_9_reset; // @[pearray.scala 209:15]
  wire  MemController_9_io_rd_valid; // @[pearray.scala 209:15]
  wire  MemController_9_io_wr_valid; // @[pearray.scala 209:15]
  wire  MemController_9_io_rd_data_valid; // @[pearray.scala 209:15]
  wire [15:0] MemController_9_io_rd_data_bits; // @[pearray.scala 209:15]
  wire  MemController_9_io_wr_data_valid; // @[pearray.scala 209:15]
  wire [15:0] MemController_9_io_wr_data_bits; // @[pearray.scala 209:15]
  wire  MemController_10_clock; // @[pearray.scala 209:15]
  wire  MemController_10_reset; // @[pearray.scala 209:15]
  wire  MemController_10_io_rd_valid; // @[pearray.scala 209:15]
  wire  MemController_10_io_wr_valid; // @[pearray.scala 209:15]
  wire  MemController_10_io_rd_data_valid; // @[pearray.scala 209:15]
  wire [15:0] MemController_10_io_rd_data_bits; // @[pearray.scala 209:15]
  wire  MemController_10_io_wr_data_valid; // @[pearray.scala 209:15]
  wire [15:0] MemController_10_io_wr_data_bits; // @[pearray.scala 209:15]
  wire  MemController_11_clock; // @[pearray.scala 209:15]
  wire  MemController_11_reset; // @[pearray.scala 209:15]
  wire  MemController_11_io_rd_valid; // @[pearray.scala 209:15]
  wire  MemController_11_io_wr_valid; // @[pearray.scala 209:15]
  wire  MemController_11_io_rd_data_valid; // @[pearray.scala 209:15]
  wire [15:0] MemController_11_io_rd_data_bits; // @[pearray.scala 209:15]
  wire  MemController_11_io_wr_data_valid; // @[pearray.scala 209:15]
  wire [15:0] MemController_11_io_wr_data_bits; // @[pearray.scala 209:15]
  wire  MemController_12_clock; // @[pearray.scala 209:15]
  wire  MemController_12_reset; // @[pearray.scala 209:15]
  wire  MemController_12_io_rd_valid; // @[pearray.scala 209:15]
  wire  MemController_12_io_wr_valid; // @[pearray.scala 209:15]
  wire  MemController_12_io_rd_data_valid; // @[pearray.scala 209:15]
  wire [15:0] MemController_12_io_rd_data_bits; // @[pearray.scala 209:15]
  wire  MemController_12_io_wr_data_valid; // @[pearray.scala 209:15]
  wire [15:0] MemController_12_io_wr_data_bits; // @[pearray.scala 209:15]
  wire  MemController_13_clock; // @[pearray.scala 209:15]
  wire  MemController_13_reset; // @[pearray.scala 209:15]
  wire  MemController_13_io_rd_valid; // @[pearray.scala 209:15]
  wire  MemController_13_io_wr_valid; // @[pearray.scala 209:15]
  wire  MemController_13_io_rd_data_valid; // @[pearray.scala 209:15]
  wire [15:0] MemController_13_io_rd_data_bits; // @[pearray.scala 209:15]
  wire  MemController_13_io_wr_data_valid; // @[pearray.scala 209:15]
  wire [15:0] MemController_13_io_wr_data_bits; // @[pearray.scala 209:15]
  wire  MemController_14_clock; // @[pearray.scala 209:15]
  wire  MemController_14_reset; // @[pearray.scala 209:15]
  wire  MemController_14_io_rd_valid; // @[pearray.scala 209:15]
  wire  MemController_14_io_wr_valid; // @[pearray.scala 209:15]
  wire  MemController_14_io_rd_data_valid; // @[pearray.scala 209:15]
  wire [15:0] MemController_14_io_rd_data_bits; // @[pearray.scala 209:15]
  wire  MemController_14_io_wr_data_valid; // @[pearray.scala 209:15]
  wire [15:0] MemController_14_io_wr_data_bits; // @[pearray.scala 209:15]
  wire  MemController_15_clock; // @[pearray.scala 209:15]
  wire  MemController_15_reset; // @[pearray.scala 209:15]
  wire  MemController_15_io_rd_valid; // @[pearray.scala 209:15]
  wire  MemController_15_io_wr_valid; // @[pearray.scala 209:15]
  wire  MemController_15_io_rd_data_valid; // @[pearray.scala 209:15]
  wire [15:0] MemController_15_io_rd_data_bits; // @[pearray.scala 209:15]
  wire  MemController_15_io_wr_data_valid; // @[pearray.scala 209:15]
  wire [15:0] MemController_15_io_wr_data_bits; // @[pearray.scala 209:15]
  wire  MemController_16_clock; // @[pearray.scala 209:15]
  wire  MemController_16_reset; // @[pearray.scala 209:15]
  wire  MemController_16_io_rd_valid; // @[pearray.scala 209:15]
  wire  MemController_16_io_wr_valid; // @[pearray.scala 209:15]
  wire  MemController_16_io_rd_data_valid; // @[pearray.scala 209:15]
  wire [15:0] MemController_16_io_rd_data_bits; // @[pearray.scala 209:15]
  wire  MemController_16_io_wr_data_valid; // @[pearray.scala 209:15]
  wire [15:0] MemController_16_io_wr_data_bits; // @[pearray.scala 209:15]
  wire  MemController_17_clock; // @[pearray.scala 209:15]
  wire  MemController_17_reset; // @[pearray.scala 209:15]
  wire  MemController_17_io_rd_valid; // @[pearray.scala 209:15]
  wire  MemController_17_io_wr_valid; // @[pearray.scala 209:15]
  wire  MemController_17_io_rd_data_valid; // @[pearray.scala 209:15]
  wire [15:0] MemController_17_io_rd_data_bits; // @[pearray.scala 209:15]
  wire  MemController_17_io_wr_data_valid; // @[pearray.scala 209:15]
  wire [15:0] MemController_17_io_wr_data_bits; // @[pearray.scala 209:15]
  wire  MemController_18_clock; // @[pearray.scala 209:15]
  wire  MemController_18_reset; // @[pearray.scala 209:15]
  wire  MemController_18_io_rd_valid; // @[pearray.scala 209:15]
  wire  MemController_18_io_wr_valid; // @[pearray.scala 209:15]
  wire  MemController_18_io_rd_data_valid; // @[pearray.scala 209:15]
  wire [15:0] MemController_18_io_rd_data_bits; // @[pearray.scala 209:15]
  wire  MemController_18_io_wr_data_valid; // @[pearray.scala 209:15]
  wire [15:0] MemController_18_io_wr_data_bits; // @[pearray.scala 209:15]
  wire  MemController_19_clock; // @[pearray.scala 209:15]
  wire  MemController_19_reset; // @[pearray.scala 209:15]
  wire  MemController_19_io_rd_valid; // @[pearray.scala 209:15]
  wire  MemController_19_io_wr_valid; // @[pearray.scala 209:15]
  wire  MemController_19_io_rd_data_valid; // @[pearray.scala 209:15]
  wire [15:0] MemController_19_io_rd_data_bits; // @[pearray.scala 209:15]
  wire  MemController_19_io_wr_data_valid; // @[pearray.scala 209:15]
  wire [15:0] MemController_19_io_wr_data_bits; // @[pearray.scala 209:15]
  wire  MemController_20_clock; // @[pearray.scala 209:15]
  wire  MemController_20_reset; // @[pearray.scala 209:15]
  wire  MemController_20_io_rd_valid; // @[pearray.scala 209:15]
  wire  MemController_20_io_wr_valid; // @[pearray.scala 209:15]
  wire  MemController_20_io_rd_data_valid; // @[pearray.scala 209:15]
  wire [15:0] MemController_20_io_rd_data_bits; // @[pearray.scala 209:15]
  wire  MemController_20_io_wr_data_valid; // @[pearray.scala 209:15]
  wire [15:0] MemController_20_io_wr_data_bits; // @[pearray.scala 209:15]
  wire  MemController_21_clock; // @[pearray.scala 209:15]
  wire  MemController_21_reset; // @[pearray.scala 209:15]
  wire  MemController_21_io_rd_valid; // @[pearray.scala 209:15]
  wire  MemController_21_io_wr_valid; // @[pearray.scala 209:15]
  wire  MemController_21_io_rd_data_valid; // @[pearray.scala 209:15]
  wire [15:0] MemController_21_io_rd_data_bits; // @[pearray.scala 209:15]
  wire  MemController_21_io_wr_data_valid; // @[pearray.scala 209:15]
  wire [15:0] MemController_21_io_wr_data_bits; // @[pearray.scala 209:15]
  wire  MemController_22_clock; // @[pearray.scala 209:15]
  wire  MemController_22_reset; // @[pearray.scala 209:15]
  wire  MemController_22_io_rd_valid; // @[pearray.scala 209:15]
  wire  MemController_22_io_wr_valid; // @[pearray.scala 209:15]
  wire  MemController_22_io_rd_data_valid; // @[pearray.scala 209:15]
  wire [15:0] MemController_22_io_rd_data_bits; // @[pearray.scala 209:15]
  wire  MemController_22_io_wr_data_valid; // @[pearray.scala 209:15]
  wire [15:0] MemController_22_io_wr_data_bits; // @[pearray.scala 209:15]
  wire  MemController_23_clock; // @[pearray.scala 209:15]
  wire  MemController_23_reset; // @[pearray.scala 209:15]
  wire  MemController_23_io_rd_valid; // @[pearray.scala 209:15]
  wire  MemController_23_io_wr_valid; // @[pearray.scala 209:15]
  wire  MemController_23_io_rd_data_valid; // @[pearray.scala 209:15]
  wire [15:0] MemController_23_io_rd_data_bits; // @[pearray.scala 209:15]
  wire  MemController_23_io_wr_data_valid; // @[pearray.scala 209:15]
  wire [15:0] MemController_23_io_wr_data_bits; // @[pearray.scala 209:15]
  wire  _T_3 = MultiDimTime_io_index_1 == 18'h0; // @[pearray.scala 182:41]
  wire  _T_4 = MultiDimTime_io_index_0 == 18'h0; // @[pearray.scala 182:89]
  wire  _T_5 = _T_3 & _T_4; // @[pearray.scala 182:67]
  reg  _T_12_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_0;
  reg  _T_12_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_1;
  reg  _T_12_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_2;
  reg  _T_12_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_3;
  wire  _T_13 = MultiDimTime_io_index_1 == 18'h1; // @[pearray.scala 182:41]
  wire  _T_15 = _T_13 & _T_4; // @[pearray.scala 182:67]
  reg  _T_22_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_4;
  reg  _T_22_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_5;
  reg  _T_22_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_6;
  reg  _T_22_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_7;
  wire  _T_23 = MultiDimTime_io_index_1 == 18'h2; // @[pearray.scala 182:41]
  wire  _T_25 = _T_23 & _T_4; // @[pearray.scala 182:67]
  reg  _T_32_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_8;
  reg  _T_32_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_9;
  reg  _T_32_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_10;
  reg  _T_32_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_11;
  wire  _T_33 = MultiDimTime_io_index_1 == 18'h3; // @[pearray.scala 182:41]
  wire  _T_35 = _T_33 & _T_4; // @[pearray.scala 182:67]
  reg  _T_42_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_12;
  reg  _T_42_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_13;
  reg  _T_42_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_14;
  reg  _T_42_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_15;
  wire  _T_43 = MultiDimTime_io_index_1 == 18'h4; // @[pearray.scala 182:41]
  wire  _T_45 = _T_43 & _T_4; // @[pearray.scala 182:67]
  reg  _T_52_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_16;
  reg  _T_52_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_17;
  reg  _T_52_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_18;
  reg  _T_52_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_19;
  wire  _T_53 = MultiDimTime_io_index_1 == 18'h5; // @[pearray.scala 182:41]
  wire  _T_55 = _T_53 & _T_4; // @[pearray.scala 182:67]
  reg  _T_62_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_20;
  reg  _T_62_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_21;
  reg  _T_62_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_22;
  reg  _T_62_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_23;
  wire  _T_63 = MultiDimTime_io_index_1 == 18'h6; // @[pearray.scala 182:41]
  wire  _T_65 = _T_63 & _T_4; // @[pearray.scala 182:67]
  reg  _T_72_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_24;
  reg  _T_72_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_25;
  reg  _T_72_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_26;
  reg  _T_72_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_27;
  wire  _T_73 = MultiDimTime_io_index_1 == 18'h7; // @[pearray.scala 182:41]
  wire  _T_75 = _T_73 & _T_4; // @[pearray.scala 182:67]
  reg  _T_82_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_28;
  reg  _T_82_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_29;
  reg  _T_82_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_30;
  reg  _T_82_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_31;
  reg  _T_92_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_32;
  reg  _T_92_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_33;
  reg  _T_92_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_34;
  reg  _T_92_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_35;
  reg  _T_102_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_36;
  reg  _T_102_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_37;
  reg  _T_102_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_38;
  reg  _T_102_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_39;
  reg  _T_112_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_40;
  reg  _T_112_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_41;
  reg  _T_112_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_42;
  reg  _T_112_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_43;
  reg  _T_122_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_44;
  reg  _T_122_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_45;
  reg  _T_122_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_46;
  reg  _T_122_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_47;
  reg  _T_132_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_48;
  reg  _T_132_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_49;
  reg  _T_132_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_50;
  reg  _T_132_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_51;
  reg  _T_142_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_52;
  reg  _T_142_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_53;
  reg  _T_142_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_54;
  reg  _T_142_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_55;
  reg  _T_152_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_56;
  reg  _T_152_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_57;
  reg  _T_152_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_58;
  reg  _T_152_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_59;
  wire  _T_153 = MultiDimTime_io_index_1 == 18'h8; // @[pearray.scala 182:41]
  wire  _T_155 = _T_153 & _T_4; // @[pearray.scala 182:67]
  reg  _T_162_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_60;
  reg  _T_162_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_61;
  reg  _T_162_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_62;
  reg  _T_162_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_63;
  reg  _T_172_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_64;
  reg  _T_172_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_65;
  reg  _T_172_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_66;
  reg  _T_172_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_67;
  reg  _T_182_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_68;
  reg  _T_182_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_69;
  reg  _T_182_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_70;
  reg  _T_182_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_71;
  reg  _T_192_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_72;
  reg  _T_192_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_73;
  reg  _T_192_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_74;
  reg  _T_192_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_75;
  reg  _T_202_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_76;
  reg  _T_202_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_77;
  reg  _T_202_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_78;
  reg  _T_202_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_79;
  reg  _T_212_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_80;
  reg  _T_212_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_81;
  reg  _T_212_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_82;
  reg  _T_212_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_83;
  reg  _T_222_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_84;
  reg  _T_222_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_85;
  reg  _T_222_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_86;
  reg  _T_222_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_87;
  reg  _T_232_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_88;
  reg  _T_232_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_89;
  reg  _T_232_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_90;
  reg  _T_232_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_91;
  wire  _T_233 = MultiDimTime_io_index_1 == 18'h9; // @[pearray.scala 182:41]
  wire  _T_235 = _T_233 & _T_4; // @[pearray.scala 182:67]
  reg  _T_242_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_92;
  reg  _T_242_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_93;
  reg  _T_242_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_94;
  reg  _T_242_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_95;
  reg  _T_252_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_96;
  reg  _T_252_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_97;
  reg  _T_252_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_98;
  reg  _T_252_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_99;
  reg  _T_262_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_100;
  reg  _T_262_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_101;
  reg  _T_262_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_102;
  reg  _T_262_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_103;
  reg  _T_272_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_104;
  reg  _T_272_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_105;
  reg  _T_272_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_106;
  reg  _T_272_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_107;
  reg  _T_282_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_108;
  reg  _T_282_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_109;
  reg  _T_282_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_110;
  reg  _T_282_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_111;
  reg  _T_292_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_112;
  reg  _T_292_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_113;
  reg  _T_292_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_114;
  reg  _T_292_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_115;
  reg  _T_302_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_116;
  reg  _T_302_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_117;
  reg  _T_302_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_118;
  reg  _T_302_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_119;
  reg  _T_312_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_120;
  reg  _T_312_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_121;
  reg  _T_312_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_122;
  reg  _T_312_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_123;
  wire  _T_313 = MultiDimTime_io_index_1 == 18'ha; // @[pearray.scala 182:41]
  wire  _T_315 = _T_313 & _T_4; // @[pearray.scala 182:67]
  reg  _T_322_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_124;
  reg  _T_322_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_125;
  reg  _T_322_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_126;
  reg  _T_322_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_127;
  reg  _T_332_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_128;
  reg  _T_332_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_129;
  reg  _T_332_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_130;
  reg  _T_332_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_131;
  reg  _T_342_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_132;
  reg  _T_342_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_133;
  reg  _T_342_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_134;
  reg  _T_342_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_135;
  reg  _T_352_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_136;
  reg  _T_352_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_137;
  reg  _T_352_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_138;
  reg  _T_352_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_139;
  reg  _T_362_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_140;
  reg  _T_362_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_141;
  reg  _T_362_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_142;
  reg  _T_362_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_143;
  reg  _T_372_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_144;
  reg  _T_372_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_145;
  reg  _T_372_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_146;
  reg  _T_372_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_147;
  reg  _T_382_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_148;
  reg  _T_382_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_149;
  reg  _T_382_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_150;
  reg  _T_382_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_151;
  reg  _T_392_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_152;
  reg  _T_392_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_153;
  reg  _T_392_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_154;
  reg  _T_392_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_155;
  wire  _T_393 = MultiDimTime_io_index_1 == 18'hb; // @[pearray.scala 182:41]
  wire  _T_395 = _T_393 & _T_4; // @[pearray.scala 182:67]
  reg  _T_402_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_156;
  reg  _T_402_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_157;
  reg  _T_402_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_158;
  reg  _T_402_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_159;
  reg  _T_412_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_160;
  reg  _T_412_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_161;
  reg  _T_412_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_162;
  reg  _T_412_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_163;
  reg  _T_422_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_164;
  reg  _T_422_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_165;
  reg  _T_422_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_166;
  reg  _T_422_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_167;
  reg  _T_432_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_168;
  reg  _T_432_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_169;
  reg  _T_432_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_170;
  reg  _T_432_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_171;
  reg  _T_442_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_172;
  reg  _T_442_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_173;
  reg  _T_442_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_174;
  reg  _T_442_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_175;
  reg  _T_452_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_176;
  reg  _T_452_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_177;
  reg  _T_452_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_178;
  reg  _T_452_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_179;
  reg  _T_462_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_180;
  reg  _T_462_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_181;
  reg  _T_462_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_182;
  reg  _T_462_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_183;
  reg  _T_472_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_184;
  reg  _T_472_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_185;
  reg  _T_472_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_186;
  reg  _T_472_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_187;
  wire  _T_473 = MultiDimTime_io_index_1 == 18'hc; // @[pearray.scala 182:41]
  wire  _T_475 = _T_473 & _T_4; // @[pearray.scala 182:67]
  reg  _T_482_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_188;
  reg  _T_482_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_189;
  reg  _T_482_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_190;
  reg  _T_482_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_191;
  reg  _T_492_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_192;
  reg  _T_492_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_193;
  reg  _T_492_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_194;
  reg  _T_492_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_195;
  reg  _T_502_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_196;
  reg  _T_502_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_197;
  reg  _T_502_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_198;
  reg  _T_502_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_199;
  reg  _T_512_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_200;
  reg  _T_512_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_201;
  reg  _T_512_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_202;
  reg  _T_512_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_203;
  reg  _T_522_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_204;
  reg  _T_522_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_205;
  reg  _T_522_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_206;
  reg  _T_522_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_207;
  reg  _T_532_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_208;
  reg  _T_532_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_209;
  reg  _T_532_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_210;
  reg  _T_532_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_211;
  reg  _T_542_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_212;
  reg  _T_542_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_213;
  reg  _T_542_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_214;
  reg  _T_542_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_215;
  reg  _T_552_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_216;
  reg  _T_552_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_217;
  reg  _T_552_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_218;
  reg  _T_552_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_219;
  wire  _T_553 = MultiDimTime_io_index_1 == 18'hd; // @[pearray.scala 182:41]
  wire  _T_555 = _T_553 & _T_4; // @[pearray.scala 182:67]
  reg  _T_562_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_220;
  reg  _T_562_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_221;
  reg  _T_562_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_222;
  reg  _T_562_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_223;
  reg  _T_572_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_224;
  reg  _T_572_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_225;
  reg  _T_572_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_226;
  reg  _T_572_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_227;
  reg  _T_582_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_228;
  reg  _T_582_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_229;
  reg  _T_582_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_230;
  reg  _T_582_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_231;
  reg  _T_592_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_232;
  reg  _T_592_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_233;
  reg  _T_592_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_234;
  reg  _T_592_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_235;
  reg  _T_602_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_236;
  reg  _T_602_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_237;
  reg  _T_602_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_238;
  reg  _T_602_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_239;
  reg  _T_612_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_240;
  reg  _T_612_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_241;
  reg  _T_612_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_242;
  reg  _T_612_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_243;
  reg  _T_622_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_244;
  reg  _T_622_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_245;
  reg  _T_622_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_246;
  reg  _T_622_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_247;
  reg  _T_632_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_248;
  reg  _T_632_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_249;
  reg  _T_632_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_250;
  reg  _T_632_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_251;
  wire  _T_633 = MultiDimTime_io_index_1 == 18'he; // @[pearray.scala 182:41]
  wire  _T_635 = _T_633 & _T_4; // @[pearray.scala 182:67]
  reg  _T_642_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_252;
  reg  _T_642_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_253;
  reg  _T_642_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_254;
  reg  _T_642_3; // @[pearray.scala 51:27]
  reg [31:0] _RAND_255;
  wire  _T_649 = MultiDimTime_io_index_1 < 18'h8; // @[pearray.scala 248:134]
  wire  _T_650 = io_exec_valid & _T_649; // @[pearray.scala 248:112]
  reg  _T_655_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_256;
  reg  _T_655_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_257;
  reg  _T_655_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_258;
  wire  _T_656 = MultiDimTime_io_index_1 >= 18'h1; // @[pearray.scala 248:82]
  wire  _T_657 = io_exec_valid & _T_656; // @[pearray.scala 248:60]
  wire  _T_658 = MultiDimTime_io_index_1 < 18'h9; // @[pearray.scala 248:134]
  wire  _T_659 = _T_657 & _T_658; // @[pearray.scala 248:112]
  reg  _T_664_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_259;
  reg  _T_664_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_260;
  reg  _T_664_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_261;
  wire  _T_665 = MultiDimTime_io_index_1 >= 18'h2; // @[pearray.scala 248:82]
  wire  _T_666 = io_exec_valid & _T_665; // @[pearray.scala 248:60]
  wire  _T_667 = MultiDimTime_io_index_1 < 18'ha; // @[pearray.scala 248:134]
  wire  _T_668 = _T_666 & _T_667; // @[pearray.scala 248:112]
  reg  _T_673_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_262;
  reg  _T_673_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_263;
  reg  _T_673_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_264;
  wire  _T_674 = MultiDimTime_io_index_1 >= 18'h3; // @[pearray.scala 248:82]
  wire  _T_675 = io_exec_valid & _T_674; // @[pearray.scala 248:60]
  wire  _T_676 = MultiDimTime_io_index_1 < 18'hb; // @[pearray.scala 248:134]
  wire  _T_677 = _T_675 & _T_676; // @[pearray.scala 248:112]
  reg  _T_682_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_265;
  reg  _T_682_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_266;
  reg  _T_682_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_267;
  wire  _T_683 = MultiDimTime_io_index_1 >= 18'h4; // @[pearray.scala 248:82]
  wire  _T_684 = io_exec_valid & _T_683; // @[pearray.scala 248:60]
  wire  _T_685 = MultiDimTime_io_index_1 < 18'hc; // @[pearray.scala 248:134]
  wire  _T_686 = _T_684 & _T_685; // @[pearray.scala 248:112]
  reg  _T_691_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_268;
  reg  _T_691_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_269;
  reg  _T_691_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_270;
  wire  _T_692 = MultiDimTime_io_index_1 >= 18'h5; // @[pearray.scala 248:82]
  wire  _T_693 = io_exec_valid & _T_692; // @[pearray.scala 248:60]
  wire  _T_694 = MultiDimTime_io_index_1 < 18'hd; // @[pearray.scala 248:134]
  wire  _T_695 = _T_693 & _T_694; // @[pearray.scala 248:112]
  reg  _T_700_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_271;
  reg  _T_700_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_272;
  reg  _T_700_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_273;
  wire  _T_701 = MultiDimTime_io_index_1 >= 18'h6; // @[pearray.scala 248:82]
  wire  _T_702 = io_exec_valid & _T_701; // @[pearray.scala 248:60]
  wire  _T_703 = MultiDimTime_io_index_1 < 18'he; // @[pearray.scala 248:134]
  wire  _T_704 = _T_702 & _T_703; // @[pearray.scala 248:112]
  reg  _T_709_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_274;
  reg  _T_709_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_275;
  reg  _T_709_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_276;
  wire  _T_710 = MultiDimTime_io_index_1 >= 18'h7; // @[pearray.scala 248:82]
  wire  _T_711 = io_exec_valid & _T_710; // @[pearray.scala 248:60]
  wire  _T_712 = MultiDimTime_io_index_1 < 18'hf; // @[pearray.scala 248:134]
  wire  _T_713 = _T_711 & _T_712; // @[pearray.scala 248:112]
  reg  _T_718_0; // @[pearray.scala 51:27]
  reg [31:0] _RAND_277;
  reg  _T_718_1; // @[pearray.scala 51:27]
  reg [31:0] _RAND_278;
  reg  _T_718_2; // @[pearray.scala 51:27]
  reg [31:0] _RAND_279;
  reg  _T_720_0; // @[pearray.scala 224:27]
  reg [31:0] _RAND_280;
  reg  _T_720_1; // @[pearray.scala 224:27]
  reg [31:0] _RAND_281;
  reg  _T_720_2; // @[pearray.scala 224:27]
  reg [31:0] _RAND_282;
  reg  _T_720_3; // @[pearray.scala 224:27]
  reg [31:0] _RAND_283;
  reg  _T_720_4; // @[pearray.scala 224:27]
  reg [31:0] _RAND_284;
  reg  _T_720_5; // @[pearray.scala 224:27]
  reg [31:0] _RAND_285;
  reg  _T_720_6; // @[pearray.scala 224:27]
  reg [31:0] _RAND_286;
  MultiDimTime MultiDimTime ( // @[pearray.scala 63:25]
    .clock(MultiDimTime_clock),
    .reset(MultiDimTime_reset),
    .io_in(MultiDimTime_io_in),
    .io_out_0(MultiDimTime_io_out_0),
    .io_out_1(MultiDimTime_io_out_1),
    .io_index_0(MultiDimTime_io_index_0),
    .io_index_1(MultiDimTime_io_index_1)
  );
  PE PE ( // @[pearray.scala 103:13]
    .clock(PE_clock),
    .reset(PE_reset),
    .io_data_2_in_valid(PE_io_data_2_in_valid),
    .io_data_2_in_bits(PE_io_data_2_in_bits),
    .io_data_2_out_valid(PE_io_data_2_out_valid),
    .io_data_2_out_bits(PE_io_data_2_out_bits),
    .io_data_1_in_valid(PE_io_data_1_in_valid),
    .io_data_1_in_bits(PE_io_data_1_in_bits),
    .io_data_1_out_valid(PE_io_data_1_out_valid),
    .io_data_1_out_bits(PE_io_data_1_out_bits),
    .io_data_0_in_valid(PE_io_data_0_in_valid),
    .io_data_0_in_bits(PE_io_data_0_in_bits),
    .io_data_0_out_valid(PE_io_data_0_out_valid),
    .io_data_0_out_bits(PE_io_data_0_out_bits),
    .io_sig_stat2trans(PE_io_sig_stat2trans)
  );
  PE PE_1 ( // @[pearray.scala 103:13]
    .clock(PE_1_clock),
    .reset(PE_1_reset),
    .io_data_2_in_valid(PE_1_io_data_2_in_valid),
    .io_data_2_in_bits(PE_1_io_data_2_in_bits),
    .io_data_2_out_valid(PE_1_io_data_2_out_valid),
    .io_data_2_out_bits(PE_1_io_data_2_out_bits),
    .io_data_1_in_valid(PE_1_io_data_1_in_valid),
    .io_data_1_in_bits(PE_1_io_data_1_in_bits),
    .io_data_1_out_valid(PE_1_io_data_1_out_valid),
    .io_data_1_out_bits(PE_1_io_data_1_out_bits),
    .io_data_0_in_valid(PE_1_io_data_0_in_valid),
    .io_data_0_in_bits(PE_1_io_data_0_in_bits),
    .io_data_0_out_valid(PE_1_io_data_0_out_valid),
    .io_data_0_out_bits(PE_1_io_data_0_out_bits),
    .io_sig_stat2trans(PE_1_io_sig_stat2trans)
  );
  PE PE_2 ( // @[pearray.scala 103:13]
    .clock(PE_2_clock),
    .reset(PE_2_reset),
    .io_data_2_in_valid(PE_2_io_data_2_in_valid),
    .io_data_2_in_bits(PE_2_io_data_2_in_bits),
    .io_data_2_out_valid(PE_2_io_data_2_out_valid),
    .io_data_2_out_bits(PE_2_io_data_2_out_bits),
    .io_data_1_in_valid(PE_2_io_data_1_in_valid),
    .io_data_1_in_bits(PE_2_io_data_1_in_bits),
    .io_data_1_out_valid(PE_2_io_data_1_out_valid),
    .io_data_1_out_bits(PE_2_io_data_1_out_bits),
    .io_data_0_in_valid(PE_2_io_data_0_in_valid),
    .io_data_0_in_bits(PE_2_io_data_0_in_bits),
    .io_data_0_out_valid(PE_2_io_data_0_out_valid),
    .io_data_0_out_bits(PE_2_io_data_0_out_bits),
    .io_sig_stat2trans(PE_2_io_sig_stat2trans)
  );
  PE PE_3 ( // @[pearray.scala 103:13]
    .clock(PE_3_clock),
    .reset(PE_3_reset),
    .io_data_2_in_valid(PE_3_io_data_2_in_valid),
    .io_data_2_in_bits(PE_3_io_data_2_in_bits),
    .io_data_2_out_valid(PE_3_io_data_2_out_valid),
    .io_data_2_out_bits(PE_3_io_data_2_out_bits),
    .io_data_1_in_valid(PE_3_io_data_1_in_valid),
    .io_data_1_in_bits(PE_3_io_data_1_in_bits),
    .io_data_1_out_valid(PE_3_io_data_1_out_valid),
    .io_data_1_out_bits(PE_3_io_data_1_out_bits),
    .io_data_0_in_valid(PE_3_io_data_0_in_valid),
    .io_data_0_in_bits(PE_3_io_data_0_in_bits),
    .io_data_0_out_valid(PE_3_io_data_0_out_valid),
    .io_data_0_out_bits(PE_3_io_data_0_out_bits),
    .io_sig_stat2trans(PE_3_io_sig_stat2trans)
  );
  PE PE_4 ( // @[pearray.scala 103:13]
    .clock(PE_4_clock),
    .reset(PE_4_reset),
    .io_data_2_in_valid(PE_4_io_data_2_in_valid),
    .io_data_2_in_bits(PE_4_io_data_2_in_bits),
    .io_data_2_out_valid(PE_4_io_data_2_out_valid),
    .io_data_2_out_bits(PE_4_io_data_2_out_bits),
    .io_data_1_in_valid(PE_4_io_data_1_in_valid),
    .io_data_1_in_bits(PE_4_io_data_1_in_bits),
    .io_data_1_out_valid(PE_4_io_data_1_out_valid),
    .io_data_1_out_bits(PE_4_io_data_1_out_bits),
    .io_data_0_in_valid(PE_4_io_data_0_in_valid),
    .io_data_0_in_bits(PE_4_io_data_0_in_bits),
    .io_data_0_out_valid(PE_4_io_data_0_out_valid),
    .io_data_0_out_bits(PE_4_io_data_0_out_bits),
    .io_sig_stat2trans(PE_4_io_sig_stat2trans)
  );
  PE PE_5 ( // @[pearray.scala 103:13]
    .clock(PE_5_clock),
    .reset(PE_5_reset),
    .io_data_2_in_valid(PE_5_io_data_2_in_valid),
    .io_data_2_in_bits(PE_5_io_data_2_in_bits),
    .io_data_2_out_valid(PE_5_io_data_2_out_valid),
    .io_data_2_out_bits(PE_5_io_data_2_out_bits),
    .io_data_1_in_valid(PE_5_io_data_1_in_valid),
    .io_data_1_in_bits(PE_5_io_data_1_in_bits),
    .io_data_1_out_valid(PE_5_io_data_1_out_valid),
    .io_data_1_out_bits(PE_5_io_data_1_out_bits),
    .io_data_0_in_valid(PE_5_io_data_0_in_valid),
    .io_data_0_in_bits(PE_5_io_data_0_in_bits),
    .io_data_0_out_valid(PE_5_io_data_0_out_valid),
    .io_data_0_out_bits(PE_5_io_data_0_out_bits),
    .io_sig_stat2trans(PE_5_io_sig_stat2trans)
  );
  PE PE_6 ( // @[pearray.scala 103:13]
    .clock(PE_6_clock),
    .reset(PE_6_reset),
    .io_data_2_in_valid(PE_6_io_data_2_in_valid),
    .io_data_2_in_bits(PE_6_io_data_2_in_bits),
    .io_data_2_out_valid(PE_6_io_data_2_out_valid),
    .io_data_2_out_bits(PE_6_io_data_2_out_bits),
    .io_data_1_in_valid(PE_6_io_data_1_in_valid),
    .io_data_1_in_bits(PE_6_io_data_1_in_bits),
    .io_data_1_out_valid(PE_6_io_data_1_out_valid),
    .io_data_1_out_bits(PE_6_io_data_1_out_bits),
    .io_data_0_in_valid(PE_6_io_data_0_in_valid),
    .io_data_0_in_bits(PE_6_io_data_0_in_bits),
    .io_data_0_out_valid(PE_6_io_data_0_out_valid),
    .io_data_0_out_bits(PE_6_io_data_0_out_bits),
    .io_sig_stat2trans(PE_6_io_sig_stat2trans)
  );
  PE PE_7 ( // @[pearray.scala 103:13]
    .clock(PE_7_clock),
    .reset(PE_7_reset),
    .io_data_2_in_valid(PE_7_io_data_2_in_valid),
    .io_data_2_in_bits(PE_7_io_data_2_in_bits),
    .io_data_2_out_valid(PE_7_io_data_2_out_valid),
    .io_data_2_out_bits(PE_7_io_data_2_out_bits),
    .io_data_1_in_valid(PE_7_io_data_1_in_valid),
    .io_data_1_in_bits(PE_7_io_data_1_in_bits),
    .io_data_1_out_valid(PE_7_io_data_1_out_valid),
    .io_data_1_out_bits(PE_7_io_data_1_out_bits),
    .io_data_0_in_valid(PE_7_io_data_0_in_valid),
    .io_data_0_in_bits(PE_7_io_data_0_in_bits),
    .io_data_0_out_valid(PE_7_io_data_0_out_valid),
    .io_data_0_out_bits(PE_7_io_data_0_out_bits),
    .io_sig_stat2trans(PE_7_io_sig_stat2trans)
  );
  PE PE_8 ( // @[pearray.scala 103:13]
    .clock(PE_8_clock),
    .reset(PE_8_reset),
    .io_data_2_in_valid(PE_8_io_data_2_in_valid),
    .io_data_2_in_bits(PE_8_io_data_2_in_bits),
    .io_data_2_out_valid(PE_8_io_data_2_out_valid),
    .io_data_2_out_bits(PE_8_io_data_2_out_bits),
    .io_data_1_in_valid(PE_8_io_data_1_in_valid),
    .io_data_1_in_bits(PE_8_io_data_1_in_bits),
    .io_data_1_out_valid(PE_8_io_data_1_out_valid),
    .io_data_1_out_bits(PE_8_io_data_1_out_bits),
    .io_data_0_in_valid(PE_8_io_data_0_in_valid),
    .io_data_0_in_bits(PE_8_io_data_0_in_bits),
    .io_data_0_out_valid(PE_8_io_data_0_out_valid),
    .io_data_0_out_bits(PE_8_io_data_0_out_bits),
    .io_sig_stat2trans(PE_8_io_sig_stat2trans)
  );
  PE PE_9 ( // @[pearray.scala 103:13]
    .clock(PE_9_clock),
    .reset(PE_9_reset),
    .io_data_2_in_valid(PE_9_io_data_2_in_valid),
    .io_data_2_in_bits(PE_9_io_data_2_in_bits),
    .io_data_2_out_valid(PE_9_io_data_2_out_valid),
    .io_data_2_out_bits(PE_9_io_data_2_out_bits),
    .io_data_1_in_valid(PE_9_io_data_1_in_valid),
    .io_data_1_in_bits(PE_9_io_data_1_in_bits),
    .io_data_1_out_valid(PE_9_io_data_1_out_valid),
    .io_data_1_out_bits(PE_9_io_data_1_out_bits),
    .io_data_0_in_valid(PE_9_io_data_0_in_valid),
    .io_data_0_in_bits(PE_9_io_data_0_in_bits),
    .io_data_0_out_valid(PE_9_io_data_0_out_valid),
    .io_data_0_out_bits(PE_9_io_data_0_out_bits),
    .io_sig_stat2trans(PE_9_io_sig_stat2trans)
  );
  PE PE_10 ( // @[pearray.scala 103:13]
    .clock(PE_10_clock),
    .reset(PE_10_reset),
    .io_data_2_in_valid(PE_10_io_data_2_in_valid),
    .io_data_2_in_bits(PE_10_io_data_2_in_bits),
    .io_data_2_out_valid(PE_10_io_data_2_out_valid),
    .io_data_2_out_bits(PE_10_io_data_2_out_bits),
    .io_data_1_in_valid(PE_10_io_data_1_in_valid),
    .io_data_1_in_bits(PE_10_io_data_1_in_bits),
    .io_data_1_out_valid(PE_10_io_data_1_out_valid),
    .io_data_1_out_bits(PE_10_io_data_1_out_bits),
    .io_data_0_in_valid(PE_10_io_data_0_in_valid),
    .io_data_0_in_bits(PE_10_io_data_0_in_bits),
    .io_data_0_out_valid(PE_10_io_data_0_out_valid),
    .io_data_0_out_bits(PE_10_io_data_0_out_bits),
    .io_sig_stat2trans(PE_10_io_sig_stat2trans)
  );
  PE PE_11 ( // @[pearray.scala 103:13]
    .clock(PE_11_clock),
    .reset(PE_11_reset),
    .io_data_2_in_valid(PE_11_io_data_2_in_valid),
    .io_data_2_in_bits(PE_11_io_data_2_in_bits),
    .io_data_2_out_valid(PE_11_io_data_2_out_valid),
    .io_data_2_out_bits(PE_11_io_data_2_out_bits),
    .io_data_1_in_valid(PE_11_io_data_1_in_valid),
    .io_data_1_in_bits(PE_11_io_data_1_in_bits),
    .io_data_1_out_valid(PE_11_io_data_1_out_valid),
    .io_data_1_out_bits(PE_11_io_data_1_out_bits),
    .io_data_0_in_valid(PE_11_io_data_0_in_valid),
    .io_data_0_in_bits(PE_11_io_data_0_in_bits),
    .io_data_0_out_valid(PE_11_io_data_0_out_valid),
    .io_data_0_out_bits(PE_11_io_data_0_out_bits),
    .io_sig_stat2trans(PE_11_io_sig_stat2trans)
  );
  PE PE_12 ( // @[pearray.scala 103:13]
    .clock(PE_12_clock),
    .reset(PE_12_reset),
    .io_data_2_in_valid(PE_12_io_data_2_in_valid),
    .io_data_2_in_bits(PE_12_io_data_2_in_bits),
    .io_data_2_out_valid(PE_12_io_data_2_out_valid),
    .io_data_2_out_bits(PE_12_io_data_2_out_bits),
    .io_data_1_in_valid(PE_12_io_data_1_in_valid),
    .io_data_1_in_bits(PE_12_io_data_1_in_bits),
    .io_data_1_out_valid(PE_12_io_data_1_out_valid),
    .io_data_1_out_bits(PE_12_io_data_1_out_bits),
    .io_data_0_in_valid(PE_12_io_data_0_in_valid),
    .io_data_0_in_bits(PE_12_io_data_0_in_bits),
    .io_data_0_out_valid(PE_12_io_data_0_out_valid),
    .io_data_0_out_bits(PE_12_io_data_0_out_bits),
    .io_sig_stat2trans(PE_12_io_sig_stat2trans)
  );
  PE PE_13 ( // @[pearray.scala 103:13]
    .clock(PE_13_clock),
    .reset(PE_13_reset),
    .io_data_2_in_valid(PE_13_io_data_2_in_valid),
    .io_data_2_in_bits(PE_13_io_data_2_in_bits),
    .io_data_2_out_valid(PE_13_io_data_2_out_valid),
    .io_data_2_out_bits(PE_13_io_data_2_out_bits),
    .io_data_1_in_valid(PE_13_io_data_1_in_valid),
    .io_data_1_in_bits(PE_13_io_data_1_in_bits),
    .io_data_1_out_valid(PE_13_io_data_1_out_valid),
    .io_data_1_out_bits(PE_13_io_data_1_out_bits),
    .io_data_0_in_valid(PE_13_io_data_0_in_valid),
    .io_data_0_in_bits(PE_13_io_data_0_in_bits),
    .io_data_0_out_valid(PE_13_io_data_0_out_valid),
    .io_data_0_out_bits(PE_13_io_data_0_out_bits),
    .io_sig_stat2trans(PE_13_io_sig_stat2trans)
  );
  PE PE_14 ( // @[pearray.scala 103:13]
    .clock(PE_14_clock),
    .reset(PE_14_reset),
    .io_data_2_in_valid(PE_14_io_data_2_in_valid),
    .io_data_2_in_bits(PE_14_io_data_2_in_bits),
    .io_data_2_out_valid(PE_14_io_data_2_out_valid),
    .io_data_2_out_bits(PE_14_io_data_2_out_bits),
    .io_data_1_in_valid(PE_14_io_data_1_in_valid),
    .io_data_1_in_bits(PE_14_io_data_1_in_bits),
    .io_data_1_out_valid(PE_14_io_data_1_out_valid),
    .io_data_1_out_bits(PE_14_io_data_1_out_bits),
    .io_data_0_in_valid(PE_14_io_data_0_in_valid),
    .io_data_0_in_bits(PE_14_io_data_0_in_bits),
    .io_data_0_out_valid(PE_14_io_data_0_out_valid),
    .io_data_0_out_bits(PE_14_io_data_0_out_bits),
    .io_sig_stat2trans(PE_14_io_sig_stat2trans)
  );
  PE PE_15 ( // @[pearray.scala 103:13]
    .clock(PE_15_clock),
    .reset(PE_15_reset),
    .io_data_2_in_valid(PE_15_io_data_2_in_valid),
    .io_data_2_in_bits(PE_15_io_data_2_in_bits),
    .io_data_2_out_valid(PE_15_io_data_2_out_valid),
    .io_data_2_out_bits(PE_15_io_data_2_out_bits),
    .io_data_1_in_valid(PE_15_io_data_1_in_valid),
    .io_data_1_in_bits(PE_15_io_data_1_in_bits),
    .io_data_1_out_valid(PE_15_io_data_1_out_valid),
    .io_data_1_out_bits(PE_15_io_data_1_out_bits),
    .io_data_0_in_valid(PE_15_io_data_0_in_valid),
    .io_data_0_in_bits(PE_15_io_data_0_in_bits),
    .io_data_0_out_valid(PE_15_io_data_0_out_valid),
    .io_data_0_out_bits(PE_15_io_data_0_out_bits),
    .io_sig_stat2trans(PE_15_io_sig_stat2trans)
  );
  PE PE_16 ( // @[pearray.scala 103:13]
    .clock(PE_16_clock),
    .reset(PE_16_reset),
    .io_data_2_in_valid(PE_16_io_data_2_in_valid),
    .io_data_2_in_bits(PE_16_io_data_2_in_bits),
    .io_data_2_out_valid(PE_16_io_data_2_out_valid),
    .io_data_2_out_bits(PE_16_io_data_2_out_bits),
    .io_data_1_in_valid(PE_16_io_data_1_in_valid),
    .io_data_1_in_bits(PE_16_io_data_1_in_bits),
    .io_data_1_out_valid(PE_16_io_data_1_out_valid),
    .io_data_1_out_bits(PE_16_io_data_1_out_bits),
    .io_data_0_in_valid(PE_16_io_data_0_in_valid),
    .io_data_0_in_bits(PE_16_io_data_0_in_bits),
    .io_data_0_out_valid(PE_16_io_data_0_out_valid),
    .io_data_0_out_bits(PE_16_io_data_0_out_bits),
    .io_sig_stat2trans(PE_16_io_sig_stat2trans)
  );
  PE PE_17 ( // @[pearray.scala 103:13]
    .clock(PE_17_clock),
    .reset(PE_17_reset),
    .io_data_2_in_valid(PE_17_io_data_2_in_valid),
    .io_data_2_in_bits(PE_17_io_data_2_in_bits),
    .io_data_2_out_valid(PE_17_io_data_2_out_valid),
    .io_data_2_out_bits(PE_17_io_data_2_out_bits),
    .io_data_1_in_valid(PE_17_io_data_1_in_valid),
    .io_data_1_in_bits(PE_17_io_data_1_in_bits),
    .io_data_1_out_valid(PE_17_io_data_1_out_valid),
    .io_data_1_out_bits(PE_17_io_data_1_out_bits),
    .io_data_0_in_valid(PE_17_io_data_0_in_valid),
    .io_data_0_in_bits(PE_17_io_data_0_in_bits),
    .io_data_0_out_valid(PE_17_io_data_0_out_valid),
    .io_data_0_out_bits(PE_17_io_data_0_out_bits),
    .io_sig_stat2trans(PE_17_io_sig_stat2trans)
  );
  PE PE_18 ( // @[pearray.scala 103:13]
    .clock(PE_18_clock),
    .reset(PE_18_reset),
    .io_data_2_in_valid(PE_18_io_data_2_in_valid),
    .io_data_2_in_bits(PE_18_io_data_2_in_bits),
    .io_data_2_out_valid(PE_18_io_data_2_out_valid),
    .io_data_2_out_bits(PE_18_io_data_2_out_bits),
    .io_data_1_in_valid(PE_18_io_data_1_in_valid),
    .io_data_1_in_bits(PE_18_io_data_1_in_bits),
    .io_data_1_out_valid(PE_18_io_data_1_out_valid),
    .io_data_1_out_bits(PE_18_io_data_1_out_bits),
    .io_data_0_in_valid(PE_18_io_data_0_in_valid),
    .io_data_0_in_bits(PE_18_io_data_0_in_bits),
    .io_data_0_out_valid(PE_18_io_data_0_out_valid),
    .io_data_0_out_bits(PE_18_io_data_0_out_bits),
    .io_sig_stat2trans(PE_18_io_sig_stat2trans)
  );
  PE PE_19 ( // @[pearray.scala 103:13]
    .clock(PE_19_clock),
    .reset(PE_19_reset),
    .io_data_2_in_valid(PE_19_io_data_2_in_valid),
    .io_data_2_in_bits(PE_19_io_data_2_in_bits),
    .io_data_2_out_valid(PE_19_io_data_2_out_valid),
    .io_data_2_out_bits(PE_19_io_data_2_out_bits),
    .io_data_1_in_valid(PE_19_io_data_1_in_valid),
    .io_data_1_in_bits(PE_19_io_data_1_in_bits),
    .io_data_1_out_valid(PE_19_io_data_1_out_valid),
    .io_data_1_out_bits(PE_19_io_data_1_out_bits),
    .io_data_0_in_valid(PE_19_io_data_0_in_valid),
    .io_data_0_in_bits(PE_19_io_data_0_in_bits),
    .io_data_0_out_valid(PE_19_io_data_0_out_valid),
    .io_data_0_out_bits(PE_19_io_data_0_out_bits),
    .io_sig_stat2trans(PE_19_io_sig_stat2trans)
  );
  PE PE_20 ( // @[pearray.scala 103:13]
    .clock(PE_20_clock),
    .reset(PE_20_reset),
    .io_data_2_in_valid(PE_20_io_data_2_in_valid),
    .io_data_2_in_bits(PE_20_io_data_2_in_bits),
    .io_data_2_out_valid(PE_20_io_data_2_out_valid),
    .io_data_2_out_bits(PE_20_io_data_2_out_bits),
    .io_data_1_in_valid(PE_20_io_data_1_in_valid),
    .io_data_1_in_bits(PE_20_io_data_1_in_bits),
    .io_data_1_out_valid(PE_20_io_data_1_out_valid),
    .io_data_1_out_bits(PE_20_io_data_1_out_bits),
    .io_data_0_in_valid(PE_20_io_data_0_in_valid),
    .io_data_0_in_bits(PE_20_io_data_0_in_bits),
    .io_data_0_out_valid(PE_20_io_data_0_out_valid),
    .io_data_0_out_bits(PE_20_io_data_0_out_bits),
    .io_sig_stat2trans(PE_20_io_sig_stat2trans)
  );
  PE PE_21 ( // @[pearray.scala 103:13]
    .clock(PE_21_clock),
    .reset(PE_21_reset),
    .io_data_2_in_valid(PE_21_io_data_2_in_valid),
    .io_data_2_in_bits(PE_21_io_data_2_in_bits),
    .io_data_2_out_valid(PE_21_io_data_2_out_valid),
    .io_data_2_out_bits(PE_21_io_data_2_out_bits),
    .io_data_1_in_valid(PE_21_io_data_1_in_valid),
    .io_data_1_in_bits(PE_21_io_data_1_in_bits),
    .io_data_1_out_valid(PE_21_io_data_1_out_valid),
    .io_data_1_out_bits(PE_21_io_data_1_out_bits),
    .io_data_0_in_valid(PE_21_io_data_0_in_valid),
    .io_data_0_in_bits(PE_21_io_data_0_in_bits),
    .io_data_0_out_valid(PE_21_io_data_0_out_valid),
    .io_data_0_out_bits(PE_21_io_data_0_out_bits),
    .io_sig_stat2trans(PE_21_io_sig_stat2trans)
  );
  PE PE_22 ( // @[pearray.scala 103:13]
    .clock(PE_22_clock),
    .reset(PE_22_reset),
    .io_data_2_in_valid(PE_22_io_data_2_in_valid),
    .io_data_2_in_bits(PE_22_io_data_2_in_bits),
    .io_data_2_out_valid(PE_22_io_data_2_out_valid),
    .io_data_2_out_bits(PE_22_io_data_2_out_bits),
    .io_data_1_in_valid(PE_22_io_data_1_in_valid),
    .io_data_1_in_bits(PE_22_io_data_1_in_bits),
    .io_data_1_out_valid(PE_22_io_data_1_out_valid),
    .io_data_1_out_bits(PE_22_io_data_1_out_bits),
    .io_data_0_in_valid(PE_22_io_data_0_in_valid),
    .io_data_0_in_bits(PE_22_io_data_0_in_bits),
    .io_data_0_out_valid(PE_22_io_data_0_out_valid),
    .io_data_0_out_bits(PE_22_io_data_0_out_bits),
    .io_sig_stat2trans(PE_22_io_sig_stat2trans)
  );
  PE PE_23 ( // @[pearray.scala 103:13]
    .clock(PE_23_clock),
    .reset(PE_23_reset),
    .io_data_2_in_valid(PE_23_io_data_2_in_valid),
    .io_data_2_in_bits(PE_23_io_data_2_in_bits),
    .io_data_2_out_valid(PE_23_io_data_2_out_valid),
    .io_data_2_out_bits(PE_23_io_data_2_out_bits),
    .io_data_1_in_valid(PE_23_io_data_1_in_valid),
    .io_data_1_in_bits(PE_23_io_data_1_in_bits),
    .io_data_1_out_valid(PE_23_io_data_1_out_valid),
    .io_data_1_out_bits(PE_23_io_data_1_out_bits),
    .io_data_0_in_valid(PE_23_io_data_0_in_valid),
    .io_data_0_in_bits(PE_23_io_data_0_in_bits),
    .io_data_0_out_valid(PE_23_io_data_0_out_valid),
    .io_data_0_out_bits(PE_23_io_data_0_out_bits),
    .io_sig_stat2trans(PE_23_io_sig_stat2trans)
  );
  PE PE_24 ( // @[pearray.scala 103:13]
    .clock(PE_24_clock),
    .reset(PE_24_reset),
    .io_data_2_in_valid(PE_24_io_data_2_in_valid),
    .io_data_2_in_bits(PE_24_io_data_2_in_bits),
    .io_data_2_out_valid(PE_24_io_data_2_out_valid),
    .io_data_2_out_bits(PE_24_io_data_2_out_bits),
    .io_data_1_in_valid(PE_24_io_data_1_in_valid),
    .io_data_1_in_bits(PE_24_io_data_1_in_bits),
    .io_data_1_out_valid(PE_24_io_data_1_out_valid),
    .io_data_1_out_bits(PE_24_io_data_1_out_bits),
    .io_data_0_in_valid(PE_24_io_data_0_in_valid),
    .io_data_0_in_bits(PE_24_io_data_0_in_bits),
    .io_data_0_out_valid(PE_24_io_data_0_out_valid),
    .io_data_0_out_bits(PE_24_io_data_0_out_bits),
    .io_sig_stat2trans(PE_24_io_sig_stat2trans)
  );
  PE PE_25 ( // @[pearray.scala 103:13]
    .clock(PE_25_clock),
    .reset(PE_25_reset),
    .io_data_2_in_valid(PE_25_io_data_2_in_valid),
    .io_data_2_in_bits(PE_25_io_data_2_in_bits),
    .io_data_2_out_valid(PE_25_io_data_2_out_valid),
    .io_data_2_out_bits(PE_25_io_data_2_out_bits),
    .io_data_1_in_valid(PE_25_io_data_1_in_valid),
    .io_data_1_in_bits(PE_25_io_data_1_in_bits),
    .io_data_1_out_valid(PE_25_io_data_1_out_valid),
    .io_data_1_out_bits(PE_25_io_data_1_out_bits),
    .io_data_0_in_valid(PE_25_io_data_0_in_valid),
    .io_data_0_in_bits(PE_25_io_data_0_in_bits),
    .io_data_0_out_valid(PE_25_io_data_0_out_valid),
    .io_data_0_out_bits(PE_25_io_data_0_out_bits),
    .io_sig_stat2trans(PE_25_io_sig_stat2trans)
  );
  PE PE_26 ( // @[pearray.scala 103:13]
    .clock(PE_26_clock),
    .reset(PE_26_reset),
    .io_data_2_in_valid(PE_26_io_data_2_in_valid),
    .io_data_2_in_bits(PE_26_io_data_2_in_bits),
    .io_data_2_out_valid(PE_26_io_data_2_out_valid),
    .io_data_2_out_bits(PE_26_io_data_2_out_bits),
    .io_data_1_in_valid(PE_26_io_data_1_in_valid),
    .io_data_1_in_bits(PE_26_io_data_1_in_bits),
    .io_data_1_out_valid(PE_26_io_data_1_out_valid),
    .io_data_1_out_bits(PE_26_io_data_1_out_bits),
    .io_data_0_in_valid(PE_26_io_data_0_in_valid),
    .io_data_0_in_bits(PE_26_io_data_0_in_bits),
    .io_data_0_out_valid(PE_26_io_data_0_out_valid),
    .io_data_0_out_bits(PE_26_io_data_0_out_bits),
    .io_sig_stat2trans(PE_26_io_sig_stat2trans)
  );
  PE PE_27 ( // @[pearray.scala 103:13]
    .clock(PE_27_clock),
    .reset(PE_27_reset),
    .io_data_2_in_valid(PE_27_io_data_2_in_valid),
    .io_data_2_in_bits(PE_27_io_data_2_in_bits),
    .io_data_2_out_valid(PE_27_io_data_2_out_valid),
    .io_data_2_out_bits(PE_27_io_data_2_out_bits),
    .io_data_1_in_valid(PE_27_io_data_1_in_valid),
    .io_data_1_in_bits(PE_27_io_data_1_in_bits),
    .io_data_1_out_valid(PE_27_io_data_1_out_valid),
    .io_data_1_out_bits(PE_27_io_data_1_out_bits),
    .io_data_0_in_valid(PE_27_io_data_0_in_valid),
    .io_data_0_in_bits(PE_27_io_data_0_in_bits),
    .io_data_0_out_valid(PE_27_io_data_0_out_valid),
    .io_data_0_out_bits(PE_27_io_data_0_out_bits),
    .io_sig_stat2trans(PE_27_io_sig_stat2trans)
  );
  PE PE_28 ( // @[pearray.scala 103:13]
    .clock(PE_28_clock),
    .reset(PE_28_reset),
    .io_data_2_in_valid(PE_28_io_data_2_in_valid),
    .io_data_2_in_bits(PE_28_io_data_2_in_bits),
    .io_data_2_out_valid(PE_28_io_data_2_out_valid),
    .io_data_2_out_bits(PE_28_io_data_2_out_bits),
    .io_data_1_in_valid(PE_28_io_data_1_in_valid),
    .io_data_1_in_bits(PE_28_io_data_1_in_bits),
    .io_data_1_out_valid(PE_28_io_data_1_out_valid),
    .io_data_1_out_bits(PE_28_io_data_1_out_bits),
    .io_data_0_in_valid(PE_28_io_data_0_in_valid),
    .io_data_0_in_bits(PE_28_io_data_0_in_bits),
    .io_data_0_out_valid(PE_28_io_data_0_out_valid),
    .io_data_0_out_bits(PE_28_io_data_0_out_bits),
    .io_sig_stat2trans(PE_28_io_sig_stat2trans)
  );
  PE PE_29 ( // @[pearray.scala 103:13]
    .clock(PE_29_clock),
    .reset(PE_29_reset),
    .io_data_2_in_valid(PE_29_io_data_2_in_valid),
    .io_data_2_in_bits(PE_29_io_data_2_in_bits),
    .io_data_2_out_valid(PE_29_io_data_2_out_valid),
    .io_data_2_out_bits(PE_29_io_data_2_out_bits),
    .io_data_1_in_valid(PE_29_io_data_1_in_valid),
    .io_data_1_in_bits(PE_29_io_data_1_in_bits),
    .io_data_1_out_valid(PE_29_io_data_1_out_valid),
    .io_data_1_out_bits(PE_29_io_data_1_out_bits),
    .io_data_0_in_valid(PE_29_io_data_0_in_valid),
    .io_data_0_in_bits(PE_29_io_data_0_in_bits),
    .io_data_0_out_valid(PE_29_io_data_0_out_valid),
    .io_data_0_out_bits(PE_29_io_data_0_out_bits),
    .io_sig_stat2trans(PE_29_io_sig_stat2trans)
  );
  PE PE_30 ( // @[pearray.scala 103:13]
    .clock(PE_30_clock),
    .reset(PE_30_reset),
    .io_data_2_in_valid(PE_30_io_data_2_in_valid),
    .io_data_2_in_bits(PE_30_io_data_2_in_bits),
    .io_data_2_out_valid(PE_30_io_data_2_out_valid),
    .io_data_2_out_bits(PE_30_io_data_2_out_bits),
    .io_data_1_in_valid(PE_30_io_data_1_in_valid),
    .io_data_1_in_bits(PE_30_io_data_1_in_bits),
    .io_data_1_out_valid(PE_30_io_data_1_out_valid),
    .io_data_1_out_bits(PE_30_io_data_1_out_bits),
    .io_data_0_in_valid(PE_30_io_data_0_in_valid),
    .io_data_0_in_bits(PE_30_io_data_0_in_bits),
    .io_data_0_out_valid(PE_30_io_data_0_out_valid),
    .io_data_0_out_bits(PE_30_io_data_0_out_bits),
    .io_sig_stat2trans(PE_30_io_sig_stat2trans)
  );
  PE PE_31 ( // @[pearray.scala 103:13]
    .clock(PE_31_clock),
    .reset(PE_31_reset),
    .io_data_2_in_valid(PE_31_io_data_2_in_valid),
    .io_data_2_in_bits(PE_31_io_data_2_in_bits),
    .io_data_2_out_valid(PE_31_io_data_2_out_valid),
    .io_data_2_out_bits(PE_31_io_data_2_out_bits),
    .io_data_1_in_valid(PE_31_io_data_1_in_valid),
    .io_data_1_in_bits(PE_31_io_data_1_in_bits),
    .io_data_1_out_valid(PE_31_io_data_1_out_valid),
    .io_data_1_out_bits(PE_31_io_data_1_out_bits),
    .io_data_0_in_valid(PE_31_io_data_0_in_valid),
    .io_data_0_in_bits(PE_31_io_data_0_in_bits),
    .io_data_0_out_valid(PE_31_io_data_0_out_valid),
    .io_data_0_out_bits(PE_31_io_data_0_out_bits),
    .io_sig_stat2trans(PE_31_io_sig_stat2trans)
  );
  PE PE_32 ( // @[pearray.scala 103:13]
    .clock(PE_32_clock),
    .reset(PE_32_reset),
    .io_data_2_in_valid(PE_32_io_data_2_in_valid),
    .io_data_2_in_bits(PE_32_io_data_2_in_bits),
    .io_data_2_out_valid(PE_32_io_data_2_out_valid),
    .io_data_2_out_bits(PE_32_io_data_2_out_bits),
    .io_data_1_in_valid(PE_32_io_data_1_in_valid),
    .io_data_1_in_bits(PE_32_io_data_1_in_bits),
    .io_data_1_out_valid(PE_32_io_data_1_out_valid),
    .io_data_1_out_bits(PE_32_io_data_1_out_bits),
    .io_data_0_in_valid(PE_32_io_data_0_in_valid),
    .io_data_0_in_bits(PE_32_io_data_0_in_bits),
    .io_data_0_out_valid(PE_32_io_data_0_out_valid),
    .io_data_0_out_bits(PE_32_io_data_0_out_bits),
    .io_sig_stat2trans(PE_32_io_sig_stat2trans)
  );
  PE PE_33 ( // @[pearray.scala 103:13]
    .clock(PE_33_clock),
    .reset(PE_33_reset),
    .io_data_2_in_valid(PE_33_io_data_2_in_valid),
    .io_data_2_in_bits(PE_33_io_data_2_in_bits),
    .io_data_2_out_valid(PE_33_io_data_2_out_valid),
    .io_data_2_out_bits(PE_33_io_data_2_out_bits),
    .io_data_1_in_valid(PE_33_io_data_1_in_valid),
    .io_data_1_in_bits(PE_33_io_data_1_in_bits),
    .io_data_1_out_valid(PE_33_io_data_1_out_valid),
    .io_data_1_out_bits(PE_33_io_data_1_out_bits),
    .io_data_0_in_valid(PE_33_io_data_0_in_valid),
    .io_data_0_in_bits(PE_33_io_data_0_in_bits),
    .io_data_0_out_valid(PE_33_io_data_0_out_valid),
    .io_data_0_out_bits(PE_33_io_data_0_out_bits),
    .io_sig_stat2trans(PE_33_io_sig_stat2trans)
  );
  PE PE_34 ( // @[pearray.scala 103:13]
    .clock(PE_34_clock),
    .reset(PE_34_reset),
    .io_data_2_in_valid(PE_34_io_data_2_in_valid),
    .io_data_2_in_bits(PE_34_io_data_2_in_bits),
    .io_data_2_out_valid(PE_34_io_data_2_out_valid),
    .io_data_2_out_bits(PE_34_io_data_2_out_bits),
    .io_data_1_in_valid(PE_34_io_data_1_in_valid),
    .io_data_1_in_bits(PE_34_io_data_1_in_bits),
    .io_data_1_out_valid(PE_34_io_data_1_out_valid),
    .io_data_1_out_bits(PE_34_io_data_1_out_bits),
    .io_data_0_in_valid(PE_34_io_data_0_in_valid),
    .io_data_0_in_bits(PE_34_io_data_0_in_bits),
    .io_data_0_out_valid(PE_34_io_data_0_out_valid),
    .io_data_0_out_bits(PE_34_io_data_0_out_bits),
    .io_sig_stat2trans(PE_34_io_sig_stat2trans)
  );
  PE PE_35 ( // @[pearray.scala 103:13]
    .clock(PE_35_clock),
    .reset(PE_35_reset),
    .io_data_2_in_valid(PE_35_io_data_2_in_valid),
    .io_data_2_in_bits(PE_35_io_data_2_in_bits),
    .io_data_2_out_valid(PE_35_io_data_2_out_valid),
    .io_data_2_out_bits(PE_35_io_data_2_out_bits),
    .io_data_1_in_valid(PE_35_io_data_1_in_valid),
    .io_data_1_in_bits(PE_35_io_data_1_in_bits),
    .io_data_1_out_valid(PE_35_io_data_1_out_valid),
    .io_data_1_out_bits(PE_35_io_data_1_out_bits),
    .io_data_0_in_valid(PE_35_io_data_0_in_valid),
    .io_data_0_in_bits(PE_35_io_data_0_in_bits),
    .io_data_0_out_valid(PE_35_io_data_0_out_valid),
    .io_data_0_out_bits(PE_35_io_data_0_out_bits),
    .io_sig_stat2trans(PE_35_io_sig_stat2trans)
  );
  PE PE_36 ( // @[pearray.scala 103:13]
    .clock(PE_36_clock),
    .reset(PE_36_reset),
    .io_data_2_in_valid(PE_36_io_data_2_in_valid),
    .io_data_2_in_bits(PE_36_io_data_2_in_bits),
    .io_data_2_out_valid(PE_36_io_data_2_out_valid),
    .io_data_2_out_bits(PE_36_io_data_2_out_bits),
    .io_data_1_in_valid(PE_36_io_data_1_in_valid),
    .io_data_1_in_bits(PE_36_io_data_1_in_bits),
    .io_data_1_out_valid(PE_36_io_data_1_out_valid),
    .io_data_1_out_bits(PE_36_io_data_1_out_bits),
    .io_data_0_in_valid(PE_36_io_data_0_in_valid),
    .io_data_0_in_bits(PE_36_io_data_0_in_bits),
    .io_data_0_out_valid(PE_36_io_data_0_out_valid),
    .io_data_0_out_bits(PE_36_io_data_0_out_bits),
    .io_sig_stat2trans(PE_36_io_sig_stat2trans)
  );
  PE PE_37 ( // @[pearray.scala 103:13]
    .clock(PE_37_clock),
    .reset(PE_37_reset),
    .io_data_2_in_valid(PE_37_io_data_2_in_valid),
    .io_data_2_in_bits(PE_37_io_data_2_in_bits),
    .io_data_2_out_valid(PE_37_io_data_2_out_valid),
    .io_data_2_out_bits(PE_37_io_data_2_out_bits),
    .io_data_1_in_valid(PE_37_io_data_1_in_valid),
    .io_data_1_in_bits(PE_37_io_data_1_in_bits),
    .io_data_1_out_valid(PE_37_io_data_1_out_valid),
    .io_data_1_out_bits(PE_37_io_data_1_out_bits),
    .io_data_0_in_valid(PE_37_io_data_0_in_valid),
    .io_data_0_in_bits(PE_37_io_data_0_in_bits),
    .io_data_0_out_valid(PE_37_io_data_0_out_valid),
    .io_data_0_out_bits(PE_37_io_data_0_out_bits),
    .io_sig_stat2trans(PE_37_io_sig_stat2trans)
  );
  PE PE_38 ( // @[pearray.scala 103:13]
    .clock(PE_38_clock),
    .reset(PE_38_reset),
    .io_data_2_in_valid(PE_38_io_data_2_in_valid),
    .io_data_2_in_bits(PE_38_io_data_2_in_bits),
    .io_data_2_out_valid(PE_38_io_data_2_out_valid),
    .io_data_2_out_bits(PE_38_io_data_2_out_bits),
    .io_data_1_in_valid(PE_38_io_data_1_in_valid),
    .io_data_1_in_bits(PE_38_io_data_1_in_bits),
    .io_data_1_out_valid(PE_38_io_data_1_out_valid),
    .io_data_1_out_bits(PE_38_io_data_1_out_bits),
    .io_data_0_in_valid(PE_38_io_data_0_in_valid),
    .io_data_0_in_bits(PE_38_io_data_0_in_bits),
    .io_data_0_out_valid(PE_38_io_data_0_out_valid),
    .io_data_0_out_bits(PE_38_io_data_0_out_bits),
    .io_sig_stat2trans(PE_38_io_sig_stat2trans)
  );
  PE PE_39 ( // @[pearray.scala 103:13]
    .clock(PE_39_clock),
    .reset(PE_39_reset),
    .io_data_2_in_valid(PE_39_io_data_2_in_valid),
    .io_data_2_in_bits(PE_39_io_data_2_in_bits),
    .io_data_2_out_valid(PE_39_io_data_2_out_valid),
    .io_data_2_out_bits(PE_39_io_data_2_out_bits),
    .io_data_1_in_valid(PE_39_io_data_1_in_valid),
    .io_data_1_in_bits(PE_39_io_data_1_in_bits),
    .io_data_1_out_valid(PE_39_io_data_1_out_valid),
    .io_data_1_out_bits(PE_39_io_data_1_out_bits),
    .io_data_0_in_valid(PE_39_io_data_0_in_valid),
    .io_data_0_in_bits(PE_39_io_data_0_in_bits),
    .io_data_0_out_valid(PE_39_io_data_0_out_valid),
    .io_data_0_out_bits(PE_39_io_data_0_out_bits),
    .io_sig_stat2trans(PE_39_io_sig_stat2trans)
  );
  PE PE_40 ( // @[pearray.scala 103:13]
    .clock(PE_40_clock),
    .reset(PE_40_reset),
    .io_data_2_in_valid(PE_40_io_data_2_in_valid),
    .io_data_2_in_bits(PE_40_io_data_2_in_bits),
    .io_data_2_out_valid(PE_40_io_data_2_out_valid),
    .io_data_2_out_bits(PE_40_io_data_2_out_bits),
    .io_data_1_in_valid(PE_40_io_data_1_in_valid),
    .io_data_1_in_bits(PE_40_io_data_1_in_bits),
    .io_data_1_out_valid(PE_40_io_data_1_out_valid),
    .io_data_1_out_bits(PE_40_io_data_1_out_bits),
    .io_data_0_in_valid(PE_40_io_data_0_in_valid),
    .io_data_0_in_bits(PE_40_io_data_0_in_bits),
    .io_data_0_out_valid(PE_40_io_data_0_out_valid),
    .io_data_0_out_bits(PE_40_io_data_0_out_bits),
    .io_sig_stat2trans(PE_40_io_sig_stat2trans)
  );
  PE PE_41 ( // @[pearray.scala 103:13]
    .clock(PE_41_clock),
    .reset(PE_41_reset),
    .io_data_2_in_valid(PE_41_io_data_2_in_valid),
    .io_data_2_in_bits(PE_41_io_data_2_in_bits),
    .io_data_2_out_valid(PE_41_io_data_2_out_valid),
    .io_data_2_out_bits(PE_41_io_data_2_out_bits),
    .io_data_1_in_valid(PE_41_io_data_1_in_valid),
    .io_data_1_in_bits(PE_41_io_data_1_in_bits),
    .io_data_1_out_valid(PE_41_io_data_1_out_valid),
    .io_data_1_out_bits(PE_41_io_data_1_out_bits),
    .io_data_0_in_valid(PE_41_io_data_0_in_valid),
    .io_data_0_in_bits(PE_41_io_data_0_in_bits),
    .io_data_0_out_valid(PE_41_io_data_0_out_valid),
    .io_data_0_out_bits(PE_41_io_data_0_out_bits),
    .io_sig_stat2trans(PE_41_io_sig_stat2trans)
  );
  PE PE_42 ( // @[pearray.scala 103:13]
    .clock(PE_42_clock),
    .reset(PE_42_reset),
    .io_data_2_in_valid(PE_42_io_data_2_in_valid),
    .io_data_2_in_bits(PE_42_io_data_2_in_bits),
    .io_data_2_out_valid(PE_42_io_data_2_out_valid),
    .io_data_2_out_bits(PE_42_io_data_2_out_bits),
    .io_data_1_in_valid(PE_42_io_data_1_in_valid),
    .io_data_1_in_bits(PE_42_io_data_1_in_bits),
    .io_data_1_out_valid(PE_42_io_data_1_out_valid),
    .io_data_1_out_bits(PE_42_io_data_1_out_bits),
    .io_data_0_in_valid(PE_42_io_data_0_in_valid),
    .io_data_0_in_bits(PE_42_io_data_0_in_bits),
    .io_data_0_out_valid(PE_42_io_data_0_out_valid),
    .io_data_0_out_bits(PE_42_io_data_0_out_bits),
    .io_sig_stat2trans(PE_42_io_sig_stat2trans)
  );
  PE PE_43 ( // @[pearray.scala 103:13]
    .clock(PE_43_clock),
    .reset(PE_43_reset),
    .io_data_2_in_valid(PE_43_io_data_2_in_valid),
    .io_data_2_in_bits(PE_43_io_data_2_in_bits),
    .io_data_2_out_valid(PE_43_io_data_2_out_valid),
    .io_data_2_out_bits(PE_43_io_data_2_out_bits),
    .io_data_1_in_valid(PE_43_io_data_1_in_valid),
    .io_data_1_in_bits(PE_43_io_data_1_in_bits),
    .io_data_1_out_valid(PE_43_io_data_1_out_valid),
    .io_data_1_out_bits(PE_43_io_data_1_out_bits),
    .io_data_0_in_valid(PE_43_io_data_0_in_valid),
    .io_data_0_in_bits(PE_43_io_data_0_in_bits),
    .io_data_0_out_valid(PE_43_io_data_0_out_valid),
    .io_data_0_out_bits(PE_43_io_data_0_out_bits),
    .io_sig_stat2trans(PE_43_io_sig_stat2trans)
  );
  PE PE_44 ( // @[pearray.scala 103:13]
    .clock(PE_44_clock),
    .reset(PE_44_reset),
    .io_data_2_in_valid(PE_44_io_data_2_in_valid),
    .io_data_2_in_bits(PE_44_io_data_2_in_bits),
    .io_data_2_out_valid(PE_44_io_data_2_out_valid),
    .io_data_2_out_bits(PE_44_io_data_2_out_bits),
    .io_data_1_in_valid(PE_44_io_data_1_in_valid),
    .io_data_1_in_bits(PE_44_io_data_1_in_bits),
    .io_data_1_out_valid(PE_44_io_data_1_out_valid),
    .io_data_1_out_bits(PE_44_io_data_1_out_bits),
    .io_data_0_in_valid(PE_44_io_data_0_in_valid),
    .io_data_0_in_bits(PE_44_io_data_0_in_bits),
    .io_data_0_out_valid(PE_44_io_data_0_out_valid),
    .io_data_0_out_bits(PE_44_io_data_0_out_bits),
    .io_sig_stat2trans(PE_44_io_sig_stat2trans)
  );
  PE PE_45 ( // @[pearray.scala 103:13]
    .clock(PE_45_clock),
    .reset(PE_45_reset),
    .io_data_2_in_valid(PE_45_io_data_2_in_valid),
    .io_data_2_in_bits(PE_45_io_data_2_in_bits),
    .io_data_2_out_valid(PE_45_io_data_2_out_valid),
    .io_data_2_out_bits(PE_45_io_data_2_out_bits),
    .io_data_1_in_valid(PE_45_io_data_1_in_valid),
    .io_data_1_in_bits(PE_45_io_data_1_in_bits),
    .io_data_1_out_valid(PE_45_io_data_1_out_valid),
    .io_data_1_out_bits(PE_45_io_data_1_out_bits),
    .io_data_0_in_valid(PE_45_io_data_0_in_valid),
    .io_data_0_in_bits(PE_45_io_data_0_in_bits),
    .io_data_0_out_valid(PE_45_io_data_0_out_valid),
    .io_data_0_out_bits(PE_45_io_data_0_out_bits),
    .io_sig_stat2trans(PE_45_io_sig_stat2trans)
  );
  PE PE_46 ( // @[pearray.scala 103:13]
    .clock(PE_46_clock),
    .reset(PE_46_reset),
    .io_data_2_in_valid(PE_46_io_data_2_in_valid),
    .io_data_2_in_bits(PE_46_io_data_2_in_bits),
    .io_data_2_out_valid(PE_46_io_data_2_out_valid),
    .io_data_2_out_bits(PE_46_io_data_2_out_bits),
    .io_data_1_in_valid(PE_46_io_data_1_in_valid),
    .io_data_1_in_bits(PE_46_io_data_1_in_bits),
    .io_data_1_out_valid(PE_46_io_data_1_out_valid),
    .io_data_1_out_bits(PE_46_io_data_1_out_bits),
    .io_data_0_in_valid(PE_46_io_data_0_in_valid),
    .io_data_0_in_bits(PE_46_io_data_0_in_bits),
    .io_data_0_out_valid(PE_46_io_data_0_out_valid),
    .io_data_0_out_bits(PE_46_io_data_0_out_bits),
    .io_sig_stat2trans(PE_46_io_sig_stat2trans)
  );
  PE PE_47 ( // @[pearray.scala 103:13]
    .clock(PE_47_clock),
    .reset(PE_47_reset),
    .io_data_2_in_valid(PE_47_io_data_2_in_valid),
    .io_data_2_in_bits(PE_47_io_data_2_in_bits),
    .io_data_2_out_valid(PE_47_io_data_2_out_valid),
    .io_data_2_out_bits(PE_47_io_data_2_out_bits),
    .io_data_1_in_valid(PE_47_io_data_1_in_valid),
    .io_data_1_in_bits(PE_47_io_data_1_in_bits),
    .io_data_1_out_valid(PE_47_io_data_1_out_valid),
    .io_data_1_out_bits(PE_47_io_data_1_out_bits),
    .io_data_0_in_valid(PE_47_io_data_0_in_valid),
    .io_data_0_in_bits(PE_47_io_data_0_in_bits),
    .io_data_0_out_valid(PE_47_io_data_0_out_valid),
    .io_data_0_out_bits(PE_47_io_data_0_out_bits),
    .io_sig_stat2trans(PE_47_io_sig_stat2trans)
  );
  PE PE_48 ( // @[pearray.scala 103:13]
    .clock(PE_48_clock),
    .reset(PE_48_reset),
    .io_data_2_in_valid(PE_48_io_data_2_in_valid),
    .io_data_2_in_bits(PE_48_io_data_2_in_bits),
    .io_data_2_out_valid(PE_48_io_data_2_out_valid),
    .io_data_2_out_bits(PE_48_io_data_2_out_bits),
    .io_data_1_in_valid(PE_48_io_data_1_in_valid),
    .io_data_1_in_bits(PE_48_io_data_1_in_bits),
    .io_data_1_out_valid(PE_48_io_data_1_out_valid),
    .io_data_1_out_bits(PE_48_io_data_1_out_bits),
    .io_data_0_in_valid(PE_48_io_data_0_in_valid),
    .io_data_0_in_bits(PE_48_io_data_0_in_bits),
    .io_data_0_out_valid(PE_48_io_data_0_out_valid),
    .io_data_0_out_bits(PE_48_io_data_0_out_bits),
    .io_sig_stat2trans(PE_48_io_sig_stat2trans)
  );
  PE PE_49 ( // @[pearray.scala 103:13]
    .clock(PE_49_clock),
    .reset(PE_49_reset),
    .io_data_2_in_valid(PE_49_io_data_2_in_valid),
    .io_data_2_in_bits(PE_49_io_data_2_in_bits),
    .io_data_2_out_valid(PE_49_io_data_2_out_valid),
    .io_data_2_out_bits(PE_49_io_data_2_out_bits),
    .io_data_1_in_valid(PE_49_io_data_1_in_valid),
    .io_data_1_in_bits(PE_49_io_data_1_in_bits),
    .io_data_1_out_valid(PE_49_io_data_1_out_valid),
    .io_data_1_out_bits(PE_49_io_data_1_out_bits),
    .io_data_0_in_valid(PE_49_io_data_0_in_valid),
    .io_data_0_in_bits(PE_49_io_data_0_in_bits),
    .io_data_0_out_valid(PE_49_io_data_0_out_valid),
    .io_data_0_out_bits(PE_49_io_data_0_out_bits),
    .io_sig_stat2trans(PE_49_io_sig_stat2trans)
  );
  PE PE_50 ( // @[pearray.scala 103:13]
    .clock(PE_50_clock),
    .reset(PE_50_reset),
    .io_data_2_in_valid(PE_50_io_data_2_in_valid),
    .io_data_2_in_bits(PE_50_io_data_2_in_bits),
    .io_data_2_out_valid(PE_50_io_data_2_out_valid),
    .io_data_2_out_bits(PE_50_io_data_2_out_bits),
    .io_data_1_in_valid(PE_50_io_data_1_in_valid),
    .io_data_1_in_bits(PE_50_io_data_1_in_bits),
    .io_data_1_out_valid(PE_50_io_data_1_out_valid),
    .io_data_1_out_bits(PE_50_io_data_1_out_bits),
    .io_data_0_in_valid(PE_50_io_data_0_in_valid),
    .io_data_0_in_bits(PE_50_io_data_0_in_bits),
    .io_data_0_out_valid(PE_50_io_data_0_out_valid),
    .io_data_0_out_bits(PE_50_io_data_0_out_bits),
    .io_sig_stat2trans(PE_50_io_sig_stat2trans)
  );
  PE PE_51 ( // @[pearray.scala 103:13]
    .clock(PE_51_clock),
    .reset(PE_51_reset),
    .io_data_2_in_valid(PE_51_io_data_2_in_valid),
    .io_data_2_in_bits(PE_51_io_data_2_in_bits),
    .io_data_2_out_valid(PE_51_io_data_2_out_valid),
    .io_data_2_out_bits(PE_51_io_data_2_out_bits),
    .io_data_1_in_valid(PE_51_io_data_1_in_valid),
    .io_data_1_in_bits(PE_51_io_data_1_in_bits),
    .io_data_1_out_valid(PE_51_io_data_1_out_valid),
    .io_data_1_out_bits(PE_51_io_data_1_out_bits),
    .io_data_0_in_valid(PE_51_io_data_0_in_valid),
    .io_data_0_in_bits(PE_51_io_data_0_in_bits),
    .io_data_0_out_valid(PE_51_io_data_0_out_valid),
    .io_data_0_out_bits(PE_51_io_data_0_out_bits),
    .io_sig_stat2trans(PE_51_io_sig_stat2trans)
  );
  PE PE_52 ( // @[pearray.scala 103:13]
    .clock(PE_52_clock),
    .reset(PE_52_reset),
    .io_data_2_in_valid(PE_52_io_data_2_in_valid),
    .io_data_2_in_bits(PE_52_io_data_2_in_bits),
    .io_data_2_out_valid(PE_52_io_data_2_out_valid),
    .io_data_2_out_bits(PE_52_io_data_2_out_bits),
    .io_data_1_in_valid(PE_52_io_data_1_in_valid),
    .io_data_1_in_bits(PE_52_io_data_1_in_bits),
    .io_data_1_out_valid(PE_52_io_data_1_out_valid),
    .io_data_1_out_bits(PE_52_io_data_1_out_bits),
    .io_data_0_in_valid(PE_52_io_data_0_in_valid),
    .io_data_0_in_bits(PE_52_io_data_0_in_bits),
    .io_data_0_out_valid(PE_52_io_data_0_out_valid),
    .io_data_0_out_bits(PE_52_io_data_0_out_bits),
    .io_sig_stat2trans(PE_52_io_sig_stat2trans)
  );
  PE PE_53 ( // @[pearray.scala 103:13]
    .clock(PE_53_clock),
    .reset(PE_53_reset),
    .io_data_2_in_valid(PE_53_io_data_2_in_valid),
    .io_data_2_in_bits(PE_53_io_data_2_in_bits),
    .io_data_2_out_valid(PE_53_io_data_2_out_valid),
    .io_data_2_out_bits(PE_53_io_data_2_out_bits),
    .io_data_1_in_valid(PE_53_io_data_1_in_valid),
    .io_data_1_in_bits(PE_53_io_data_1_in_bits),
    .io_data_1_out_valid(PE_53_io_data_1_out_valid),
    .io_data_1_out_bits(PE_53_io_data_1_out_bits),
    .io_data_0_in_valid(PE_53_io_data_0_in_valid),
    .io_data_0_in_bits(PE_53_io_data_0_in_bits),
    .io_data_0_out_valid(PE_53_io_data_0_out_valid),
    .io_data_0_out_bits(PE_53_io_data_0_out_bits),
    .io_sig_stat2trans(PE_53_io_sig_stat2trans)
  );
  PE PE_54 ( // @[pearray.scala 103:13]
    .clock(PE_54_clock),
    .reset(PE_54_reset),
    .io_data_2_in_valid(PE_54_io_data_2_in_valid),
    .io_data_2_in_bits(PE_54_io_data_2_in_bits),
    .io_data_2_out_valid(PE_54_io_data_2_out_valid),
    .io_data_2_out_bits(PE_54_io_data_2_out_bits),
    .io_data_1_in_valid(PE_54_io_data_1_in_valid),
    .io_data_1_in_bits(PE_54_io_data_1_in_bits),
    .io_data_1_out_valid(PE_54_io_data_1_out_valid),
    .io_data_1_out_bits(PE_54_io_data_1_out_bits),
    .io_data_0_in_valid(PE_54_io_data_0_in_valid),
    .io_data_0_in_bits(PE_54_io_data_0_in_bits),
    .io_data_0_out_valid(PE_54_io_data_0_out_valid),
    .io_data_0_out_bits(PE_54_io_data_0_out_bits),
    .io_sig_stat2trans(PE_54_io_sig_stat2trans)
  );
  PE PE_55 ( // @[pearray.scala 103:13]
    .clock(PE_55_clock),
    .reset(PE_55_reset),
    .io_data_2_in_valid(PE_55_io_data_2_in_valid),
    .io_data_2_in_bits(PE_55_io_data_2_in_bits),
    .io_data_2_out_valid(PE_55_io_data_2_out_valid),
    .io_data_2_out_bits(PE_55_io_data_2_out_bits),
    .io_data_1_in_valid(PE_55_io_data_1_in_valid),
    .io_data_1_in_bits(PE_55_io_data_1_in_bits),
    .io_data_1_out_valid(PE_55_io_data_1_out_valid),
    .io_data_1_out_bits(PE_55_io_data_1_out_bits),
    .io_data_0_in_valid(PE_55_io_data_0_in_valid),
    .io_data_0_in_bits(PE_55_io_data_0_in_bits),
    .io_data_0_out_valid(PE_55_io_data_0_out_valid),
    .io_data_0_out_bits(PE_55_io_data_0_out_bits),
    .io_sig_stat2trans(PE_55_io_sig_stat2trans)
  );
  PE PE_56 ( // @[pearray.scala 103:13]
    .clock(PE_56_clock),
    .reset(PE_56_reset),
    .io_data_2_in_valid(PE_56_io_data_2_in_valid),
    .io_data_2_in_bits(PE_56_io_data_2_in_bits),
    .io_data_2_out_valid(PE_56_io_data_2_out_valid),
    .io_data_2_out_bits(PE_56_io_data_2_out_bits),
    .io_data_1_in_valid(PE_56_io_data_1_in_valid),
    .io_data_1_in_bits(PE_56_io_data_1_in_bits),
    .io_data_1_out_valid(PE_56_io_data_1_out_valid),
    .io_data_1_out_bits(PE_56_io_data_1_out_bits),
    .io_data_0_in_valid(PE_56_io_data_0_in_valid),
    .io_data_0_in_bits(PE_56_io_data_0_in_bits),
    .io_data_0_out_valid(PE_56_io_data_0_out_valid),
    .io_data_0_out_bits(PE_56_io_data_0_out_bits),
    .io_sig_stat2trans(PE_56_io_sig_stat2trans)
  );
  PE PE_57 ( // @[pearray.scala 103:13]
    .clock(PE_57_clock),
    .reset(PE_57_reset),
    .io_data_2_in_valid(PE_57_io_data_2_in_valid),
    .io_data_2_in_bits(PE_57_io_data_2_in_bits),
    .io_data_2_out_valid(PE_57_io_data_2_out_valid),
    .io_data_2_out_bits(PE_57_io_data_2_out_bits),
    .io_data_1_in_valid(PE_57_io_data_1_in_valid),
    .io_data_1_in_bits(PE_57_io_data_1_in_bits),
    .io_data_1_out_valid(PE_57_io_data_1_out_valid),
    .io_data_1_out_bits(PE_57_io_data_1_out_bits),
    .io_data_0_in_valid(PE_57_io_data_0_in_valid),
    .io_data_0_in_bits(PE_57_io_data_0_in_bits),
    .io_data_0_out_valid(PE_57_io_data_0_out_valid),
    .io_data_0_out_bits(PE_57_io_data_0_out_bits),
    .io_sig_stat2trans(PE_57_io_sig_stat2trans)
  );
  PE PE_58 ( // @[pearray.scala 103:13]
    .clock(PE_58_clock),
    .reset(PE_58_reset),
    .io_data_2_in_valid(PE_58_io_data_2_in_valid),
    .io_data_2_in_bits(PE_58_io_data_2_in_bits),
    .io_data_2_out_valid(PE_58_io_data_2_out_valid),
    .io_data_2_out_bits(PE_58_io_data_2_out_bits),
    .io_data_1_in_valid(PE_58_io_data_1_in_valid),
    .io_data_1_in_bits(PE_58_io_data_1_in_bits),
    .io_data_1_out_valid(PE_58_io_data_1_out_valid),
    .io_data_1_out_bits(PE_58_io_data_1_out_bits),
    .io_data_0_in_valid(PE_58_io_data_0_in_valid),
    .io_data_0_in_bits(PE_58_io_data_0_in_bits),
    .io_data_0_out_valid(PE_58_io_data_0_out_valid),
    .io_data_0_out_bits(PE_58_io_data_0_out_bits),
    .io_sig_stat2trans(PE_58_io_sig_stat2trans)
  );
  PE PE_59 ( // @[pearray.scala 103:13]
    .clock(PE_59_clock),
    .reset(PE_59_reset),
    .io_data_2_in_valid(PE_59_io_data_2_in_valid),
    .io_data_2_in_bits(PE_59_io_data_2_in_bits),
    .io_data_2_out_valid(PE_59_io_data_2_out_valid),
    .io_data_2_out_bits(PE_59_io_data_2_out_bits),
    .io_data_1_in_valid(PE_59_io_data_1_in_valid),
    .io_data_1_in_bits(PE_59_io_data_1_in_bits),
    .io_data_1_out_valid(PE_59_io_data_1_out_valid),
    .io_data_1_out_bits(PE_59_io_data_1_out_bits),
    .io_data_0_in_valid(PE_59_io_data_0_in_valid),
    .io_data_0_in_bits(PE_59_io_data_0_in_bits),
    .io_data_0_out_valid(PE_59_io_data_0_out_valid),
    .io_data_0_out_bits(PE_59_io_data_0_out_bits),
    .io_sig_stat2trans(PE_59_io_sig_stat2trans)
  );
  PE PE_60 ( // @[pearray.scala 103:13]
    .clock(PE_60_clock),
    .reset(PE_60_reset),
    .io_data_2_in_valid(PE_60_io_data_2_in_valid),
    .io_data_2_in_bits(PE_60_io_data_2_in_bits),
    .io_data_2_out_valid(PE_60_io_data_2_out_valid),
    .io_data_2_out_bits(PE_60_io_data_2_out_bits),
    .io_data_1_in_valid(PE_60_io_data_1_in_valid),
    .io_data_1_in_bits(PE_60_io_data_1_in_bits),
    .io_data_1_out_valid(PE_60_io_data_1_out_valid),
    .io_data_1_out_bits(PE_60_io_data_1_out_bits),
    .io_data_0_in_valid(PE_60_io_data_0_in_valid),
    .io_data_0_in_bits(PE_60_io_data_0_in_bits),
    .io_data_0_out_valid(PE_60_io_data_0_out_valid),
    .io_data_0_out_bits(PE_60_io_data_0_out_bits),
    .io_sig_stat2trans(PE_60_io_sig_stat2trans)
  );
  PE PE_61 ( // @[pearray.scala 103:13]
    .clock(PE_61_clock),
    .reset(PE_61_reset),
    .io_data_2_in_valid(PE_61_io_data_2_in_valid),
    .io_data_2_in_bits(PE_61_io_data_2_in_bits),
    .io_data_2_out_valid(PE_61_io_data_2_out_valid),
    .io_data_2_out_bits(PE_61_io_data_2_out_bits),
    .io_data_1_in_valid(PE_61_io_data_1_in_valid),
    .io_data_1_in_bits(PE_61_io_data_1_in_bits),
    .io_data_1_out_valid(PE_61_io_data_1_out_valid),
    .io_data_1_out_bits(PE_61_io_data_1_out_bits),
    .io_data_0_in_valid(PE_61_io_data_0_in_valid),
    .io_data_0_in_bits(PE_61_io_data_0_in_bits),
    .io_data_0_out_valid(PE_61_io_data_0_out_valid),
    .io_data_0_out_bits(PE_61_io_data_0_out_bits),
    .io_sig_stat2trans(PE_61_io_sig_stat2trans)
  );
  PE PE_62 ( // @[pearray.scala 103:13]
    .clock(PE_62_clock),
    .reset(PE_62_reset),
    .io_data_2_in_valid(PE_62_io_data_2_in_valid),
    .io_data_2_in_bits(PE_62_io_data_2_in_bits),
    .io_data_2_out_valid(PE_62_io_data_2_out_valid),
    .io_data_2_out_bits(PE_62_io_data_2_out_bits),
    .io_data_1_in_valid(PE_62_io_data_1_in_valid),
    .io_data_1_in_bits(PE_62_io_data_1_in_bits),
    .io_data_1_out_valid(PE_62_io_data_1_out_valid),
    .io_data_1_out_bits(PE_62_io_data_1_out_bits),
    .io_data_0_in_valid(PE_62_io_data_0_in_valid),
    .io_data_0_in_bits(PE_62_io_data_0_in_bits),
    .io_data_0_out_valid(PE_62_io_data_0_out_valid),
    .io_data_0_out_bits(PE_62_io_data_0_out_bits),
    .io_sig_stat2trans(PE_62_io_sig_stat2trans)
  );
  PE PE_63 ( // @[pearray.scala 103:13]
    .clock(PE_63_clock),
    .reset(PE_63_reset),
    .io_data_2_in_valid(PE_63_io_data_2_in_valid),
    .io_data_2_in_bits(PE_63_io_data_2_in_bits),
    .io_data_2_out_valid(PE_63_io_data_2_out_valid),
    .io_data_2_out_bits(PE_63_io_data_2_out_bits),
    .io_data_1_in_valid(PE_63_io_data_1_in_valid),
    .io_data_1_in_bits(PE_63_io_data_1_in_bits),
    .io_data_1_out_valid(PE_63_io_data_1_out_valid),
    .io_data_1_out_bits(PE_63_io_data_1_out_bits),
    .io_data_0_in_valid(PE_63_io_data_0_in_valid),
    .io_data_0_in_bits(PE_63_io_data_0_in_bits),
    .io_data_0_out_valid(PE_63_io_data_0_out_valid),
    .io_data_0_out_bits(PE_63_io_data_0_out_bits),
    .io_sig_stat2trans(PE_63_io_sig_stat2trans)
  );
  PENetwork PENetwork ( // @[pearray.scala 137:13]
    .io_to_pes_0_out_valid(PENetwork_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_io_to_pes_7_out_bits),
    .io_to_mem_valid(PENetwork_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_io_to_mem_bits)
  );
  PENetwork PENetwork_1 ( // @[pearray.scala 137:13]
    .io_to_pes_0_out_valid(PENetwork_1_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_1_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_1_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_1_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_1_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_1_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_1_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_1_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_1_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_1_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_1_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_1_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_1_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_1_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_1_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_1_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_1_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_1_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_1_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_1_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_1_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_1_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_1_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_1_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_1_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_1_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_1_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_1_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_1_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_1_io_to_pes_7_out_bits),
    .io_to_mem_valid(PENetwork_1_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_1_io_to_mem_bits)
  );
  PENetwork PENetwork_2 ( // @[pearray.scala 137:13]
    .io_to_pes_0_out_valid(PENetwork_2_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_2_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_2_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_2_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_2_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_2_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_2_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_2_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_2_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_2_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_2_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_2_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_2_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_2_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_2_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_2_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_2_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_2_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_2_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_2_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_2_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_2_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_2_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_2_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_2_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_2_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_2_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_2_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_2_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_2_io_to_pes_7_out_bits),
    .io_to_mem_valid(PENetwork_2_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_2_io_to_mem_bits)
  );
  PENetwork PENetwork_3 ( // @[pearray.scala 137:13]
    .io_to_pes_0_out_valid(PENetwork_3_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_3_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_3_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_3_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_3_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_3_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_3_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_3_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_3_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_3_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_3_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_3_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_3_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_3_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_3_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_3_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_3_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_3_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_3_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_3_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_3_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_3_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_3_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_3_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_3_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_3_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_3_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_3_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_3_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_3_io_to_pes_7_out_bits),
    .io_to_mem_valid(PENetwork_3_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_3_io_to_mem_bits)
  );
  PENetwork PENetwork_4 ( // @[pearray.scala 137:13]
    .io_to_pes_0_out_valid(PENetwork_4_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_4_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_4_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_4_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_4_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_4_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_4_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_4_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_4_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_4_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_4_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_4_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_4_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_4_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_4_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_4_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_4_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_4_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_4_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_4_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_4_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_4_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_4_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_4_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_4_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_4_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_4_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_4_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_4_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_4_io_to_pes_7_out_bits),
    .io_to_mem_valid(PENetwork_4_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_4_io_to_mem_bits)
  );
  PENetwork PENetwork_5 ( // @[pearray.scala 137:13]
    .io_to_pes_0_out_valid(PENetwork_5_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_5_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_5_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_5_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_5_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_5_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_5_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_5_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_5_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_5_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_5_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_5_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_5_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_5_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_5_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_5_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_5_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_5_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_5_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_5_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_5_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_5_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_5_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_5_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_5_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_5_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_5_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_5_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_5_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_5_io_to_pes_7_out_bits),
    .io_to_mem_valid(PENetwork_5_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_5_io_to_mem_bits)
  );
  PENetwork PENetwork_6 ( // @[pearray.scala 137:13]
    .io_to_pes_0_out_valid(PENetwork_6_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_6_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_6_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_6_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_6_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_6_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_6_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_6_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_6_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_6_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_6_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_6_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_6_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_6_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_6_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_6_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_6_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_6_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_6_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_6_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_6_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_6_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_6_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_6_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_6_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_6_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_6_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_6_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_6_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_6_io_to_pes_7_out_bits),
    .io_to_mem_valid(PENetwork_6_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_6_io_to_mem_bits)
  );
  PENetwork PENetwork_7 ( // @[pearray.scala 137:13]
    .io_to_pes_0_out_valid(PENetwork_7_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_7_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_7_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_7_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_7_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_7_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_7_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_7_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_7_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_7_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_7_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_7_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_7_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_7_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_7_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_7_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_7_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_7_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_7_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_7_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_7_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_7_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_7_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_7_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_7_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_7_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_7_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_7_io_to_pes_7_in_bits),
    .io_to_pes_7_out_valid(PENetwork_7_io_to_pes_7_out_valid),
    .io_to_pes_7_out_bits(PENetwork_7_io_to_pes_7_out_bits),
    .io_to_mem_valid(PENetwork_7_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_7_io_to_mem_bits)
  );
  PENetwork_8 PENetwork_8 ( // @[pearray.scala 137:13]
    .io_to_pes_0_in_valid(PENetwork_8_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_8_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_8_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_8_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_8_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_8_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_8_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_8_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_8_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_8_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_8_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_8_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_8_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_8_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_8_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_8_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_8_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_8_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_8_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_8_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_8_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_8_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_8_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_8_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_8_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_8_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_8_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_8_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_8_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_8_io_to_pes_7_in_bits),
    .io_to_mem_valid(PENetwork_8_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_8_io_to_mem_bits)
  );
  PENetwork_8 PENetwork_9 ( // @[pearray.scala 137:13]
    .io_to_pes_0_in_valid(PENetwork_9_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_9_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_9_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_9_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_9_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_9_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_9_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_9_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_9_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_9_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_9_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_9_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_9_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_9_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_9_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_9_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_9_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_9_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_9_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_9_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_9_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_9_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_9_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_9_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_9_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_9_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_9_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_9_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_9_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_9_io_to_pes_7_in_bits),
    .io_to_mem_valid(PENetwork_9_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_9_io_to_mem_bits)
  );
  PENetwork_8 PENetwork_10 ( // @[pearray.scala 137:13]
    .io_to_pes_0_in_valid(PENetwork_10_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_10_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_10_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_10_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_10_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_10_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_10_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_10_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_10_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_10_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_10_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_10_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_10_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_10_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_10_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_10_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_10_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_10_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_10_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_10_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_10_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_10_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_10_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_10_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_10_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_10_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_10_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_10_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_10_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_10_io_to_pes_7_in_bits),
    .io_to_mem_valid(PENetwork_10_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_10_io_to_mem_bits)
  );
  PENetwork_8 PENetwork_11 ( // @[pearray.scala 137:13]
    .io_to_pes_0_in_valid(PENetwork_11_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_11_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_11_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_11_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_11_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_11_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_11_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_11_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_11_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_11_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_11_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_11_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_11_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_11_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_11_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_11_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_11_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_11_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_11_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_11_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_11_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_11_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_11_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_11_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_11_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_11_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_11_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_11_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_11_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_11_io_to_pes_7_in_bits),
    .io_to_mem_valid(PENetwork_11_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_11_io_to_mem_bits)
  );
  PENetwork_8 PENetwork_12 ( // @[pearray.scala 137:13]
    .io_to_pes_0_in_valid(PENetwork_12_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_12_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_12_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_12_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_12_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_12_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_12_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_12_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_12_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_12_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_12_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_12_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_12_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_12_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_12_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_12_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_12_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_12_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_12_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_12_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_12_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_12_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_12_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_12_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_12_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_12_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_12_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_12_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_12_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_12_io_to_pes_7_in_bits),
    .io_to_mem_valid(PENetwork_12_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_12_io_to_mem_bits)
  );
  PENetwork_8 PENetwork_13 ( // @[pearray.scala 137:13]
    .io_to_pes_0_in_valid(PENetwork_13_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_13_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_13_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_13_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_13_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_13_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_13_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_13_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_13_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_13_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_13_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_13_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_13_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_13_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_13_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_13_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_13_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_13_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_13_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_13_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_13_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_13_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_13_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_13_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_13_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_13_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_13_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_13_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_13_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_13_io_to_pes_7_in_bits),
    .io_to_mem_valid(PENetwork_13_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_13_io_to_mem_bits)
  );
  PENetwork_8 PENetwork_14 ( // @[pearray.scala 137:13]
    .io_to_pes_0_in_valid(PENetwork_14_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_14_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_14_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_14_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_14_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_14_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_14_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_14_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_14_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_14_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_14_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_14_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_14_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_14_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_14_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_14_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_14_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_14_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_14_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_14_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_14_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_14_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_14_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_14_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_14_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_14_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_14_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_14_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_14_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_14_io_to_pes_7_in_bits),
    .io_to_mem_valid(PENetwork_14_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_14_io_to_mem_bits)
  );
  PENetwork_8 PENetwork_15 ( // @[pearray.scala 137:13]
    .io_to_pes_0_in_valid(PENetwork_15_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_15_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_15_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_15_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_15_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_15_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_15_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_15_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_15_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_15_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_15_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_15_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_15_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_15_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_15_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_15_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_15_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_15_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_15_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_15_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_15_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_15_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_15_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_15_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_15_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_15_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_15_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_15_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_15_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_15_io_to_pes_7_in_bits),
    .io_to_mem_valid(PENetwork_15_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_15_io_to_mem_bits)
  );
  PENetwork_8 PENetwork_16 ( // @[pearray.scala 137:13]
    .io_to_pes_0_in_valid(PENetwork_16_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_16_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_16_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_16_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_16_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_16_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_16_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_16_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_16_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_16_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_16_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_16_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_16_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_16_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_16_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_16_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_16_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_16_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_16_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_16_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_16_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_16_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_16_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_16_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_16_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_16_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_16_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_16_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_16_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_16_io_to_pes_7_in_bits),
    .io_to_mem_valid(PENetwork_16_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_16_io_to_mem_bits)
  );
  PENetwork_8 PENetwork_17 ( // @[pearray.scala 137:13]
    .io_to_pes_0_in_valid(PENetwork_17_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_17_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_17_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_17_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_17_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_17_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_17_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_17_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_17_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_17_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_17_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_17_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_17_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_17_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_17_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_17_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_17_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_17_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_17_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_17_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_17_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_17_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_17_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_17_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_17_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_17_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_17_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_17_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_17_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_17_io_to_pes_7_in_bits),
    .io_to_mem_valid(PENetwork_17_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_17_io_to_mem_bits)
  );
  PENetwork_8 PENetwork_18 ( // @[pearray.scala 137:13]
    .io_to_pes_0_in_valid(PENetwork_18_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_18_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_18_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_18_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_18_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_18_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_18_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_18_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_18_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_18_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_18_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_18_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_18_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_18_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_18_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_18_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_18_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_18_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_18_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_18_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_18_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_18_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_18_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_18_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_18_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_18_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_18_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_18_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_18_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_18_io_to_pes_7_in_bits),
    .io_to_mem_valid(PENetwork_18_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_18_io_to_mem_bits)
  );
  PENetwork_8 PENetwork_19 ( // @[pearray.scala 137:13]
    .io_to_pes_0_in_valid(PENetwork_19_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_19_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_19_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_19_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_19_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_19_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_19_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_19_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_19_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_19_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_19_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_19_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_19_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_19_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_19_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_19_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_19_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_19_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_19_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_19_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_19_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_19_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_19_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_19_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_19_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_19_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_19_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_19_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_19_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_19_io_to_pes_7_in_bits),
    .io_to_mem_valid(PENetwork_19_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_19_io_to_mem_bits)
  );
  PENetwork_8 PENetwork_20 ( // @[pearray.scala 137:13]
    .io_to_pes_0_in_valid(PENetwork_20_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_20_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_20_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_20_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_20_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_20_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_20_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_20_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_20_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_20_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_20_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_20_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_20_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_20_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_20_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_20_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_20_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_20_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_20_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_20_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_20_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_20_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_20_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_20_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_20_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_20_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_20_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_20_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_20_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_20_io_to_pes_7_in_bits),
    .io_to_mem_valid(PENetwork_20_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_20_io_to_mem_bits)
  );
  PENetwork_8 PENetwork_21 ( // @[pearray.scala 137:13]
    .io_to_pes_0_in_valid(PENetwork_21_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_21_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_21_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_21_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_21_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_21_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_21_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_21_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_21_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_21_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_21_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_21_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_21_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_21_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_21_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_21_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_21_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_21_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_21_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_21_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_21_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_21_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_21_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_21_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_21_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_21_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_21_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_21_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_21_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_21_io_to_pes_7_in_bits),
    .io_to_mem_valid(PENetwork_21_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_21_io_to_mem_bits)
  );
  PENetwork_8 PENetwork_22 ( // @[pearray.scala 137:13]
    .io_to_pes_0_in_valid(PENetwork_22_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_22_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_22_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_22_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_22_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_22_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_22_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_22_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_22_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_22_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_22_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_22_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_22_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_22_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_22_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_22_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_22_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_22_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_22_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_22_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_22_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_22_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_22_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_22_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_22_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_22_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_22_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_22_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_22_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_22_io_to_pes_7_in_bits),
    .io_to_mem_valid(PENetwork_22_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_22_io_to_mem_bits)
  );
  PENetwork_8 PENetwork_23 ( // @[pearray.scala 137:13]
    .io_to_pes_0_in_valid(PENetwork_23_io_to_pes_0_in_valid),
    .io_to_pes_0_in_bits(PENetwork_23_io_to_pes_0_in_bits),
    .io_to_pes_0_out_valid(PENetwork_23_io_to_pes_0_out_valid),
    .io_to_pes_0_out_bits(PENetwork_23_io_to_pes_0_out_bits),
    .io_to_pes_1_in_valid(PENetwork_23_io_to_pes_1_in_valid),
    .io_to_pes_1_in_bits(PENetwork_23_io_to_pes_1_in_bits),
    .io_to_pes_1_out_valid(PENetwork_23_io_to_pes_1_out_valid),
    .io_to_pes_1_out_bits(PENetwork_23_io_to_pes_1_out_bits),
    .io_to_pes_2_in_valid(PENetwork_23_io_to_pes_2_in_valid),
    .io_to_pes_2_in_bits(PENetwork_23_io_to_pes_2_in_bits),
    .io_to_pes_2_out_valid(PENetwork_23_io_to_pes_2_out_valid),
    .io_to_pes_2_out_bits(PENetwork_23_io_to_pes_2_out_bits),
    .io_to_pes_3_in_valid(PENetwork_23_io_to_pes_3_in_valid),
    .io_to_pes_3_in_bits(PENetwork_23_io_to_pes_3_in_bits),
    .io_to_pes_3_out_valid(PENetwork_23_io_to_pes_3_out_valid),
    .io_to_pes_3_out_bits(PENetwork_23_io_to_pes_3_out_bits),
    .io_to_pes_4_in_valid(PENetwork_23_io_to_pes_4_in_valid),
    .io_to_pes_4_in_bits(PENetwork_23_io_to_pes_4_in_bits),
    .io_to_pes_4_out_valid(PENetwork_23_io_to_pes_4_out_valid),
    .io_to_pes_4_out_bits(PENetwork_23_io_to_pes_4_out_bits),
    .io_to_pes_5_in_valid(PENetwork_23_io_to_pes_5_in_valid),
    .io_to_pes_5_in_bits(PENetwork_23_io_to_pes_5_in_bits),
    .io_to_pes_5_out_valid(PENetwork_23_io_to_pes_5_out_valid),
    .io_to_pes_5_out_bits(PENetwork_23_io_to_pes_5_out_bits),
    .io_to_pes_6_in_valid(PENetwork_23_io_to_pes_6_in_valid),
    .io_to_pes_6_in_bits(PENetwork_23_io_to_pes_6_in_bits),
    .io_to_pes_6_out_valid(PENetwork_23_io_to_pes_6_out_valid),
    .io_to_pes_6_out_bits(PENetwork_23_io_to_pes_6_out_bits),
    .io_to_pes_7_in_valid(PENetwork_23_io_to_pes_7_in_valid),
    .io_to_pes_7_in_bits(PENetwork_23_io_to_pes_7_in_bits),
    .io_to_mem_valid(PENetwork_23_io_to_mem_valid),
    .io_to_mem_bits(PENetwork_23_io_to_mem_bits)
  );
  MemController MemController ( // @[pearray.scala 211:15]
    .clock(MemController_clock),
    .reset(MemController_reset),
    .io_rd_valid(MemController_io_rd_valid),
    .io_wr_valid(MemController_io_wr_valid),
    .io_rd_data_valid(MemController_io_rd_data_valid),
    .io_rd_data_bits(MemController_io_rd_data_bits),
    .io_wr_data_valid(MemController_io_wr_data_valid),
    .io_wr_data_bits(MemController_io_wr_data_bits)
  );
  MemController MemController_1 ( // @[pearray.scala 211:15]
    .clock(MemController_1_clock),
    .reset(MemController_1_reset),
    .io_rd_valid(MemController_1_io_rd_valid),
    .io_wr_valid(MemController_1_io_wr_valid),
    .io_rd_data_valid(MemController_1_io_rd_data_valid),
    .io_rd_data_bits(MemController_1_io_rd_data_bits),
    .io_wr_data_valid(MemController_1_io_wr_data_valid),
    .io_wr_data_bits(MemController_1_io_wr_data_bits)
  );
  MemController MemController_2 ( // @[pearray.scala 211:15]
    .clock(MemController_2_clock),
    .reset(MemController_2_reset),
    .io_rd_valid(MemController_2_io_rd_valid),
    .io_wr_valid(MemController_2_io_wr_valid),
    .io_rd_data_valid(MemController_2_io_rd_data_valid),
    .io_rd_data_bits(MemController_2_io_rd_data_bits),
    .io_wr_data_valid(MemController_2_io_wr_data_valid),
    .io_wr_data_bits(MemController_2_io_wr_data_bits)
  );
  MemController MemController_3 ( // @[pearray.scala 211:15]
    .clock(MemController_3_clock),
    .reset(MemController_3_reset),
    .io_rd_valid(MemController_3_io_rd_valid),
    .io_wr_valid(MemController_3_io_wr_valid),
    .io_rd_data_valid(MemController_3_io_rd_data_valid),
    .io_rd_data_bits(MemController_3_io_rd_data_bits),
    .io_wr_data_valid(MemController_3_io_wr_data_valid),
    .io_wr_data_bits(MemController_3_io_wr_data_bits)
  );
  MemController MemController_4 ( // @[pearray.scala 211:15]
    .clock(MemController_4_clock),
    .reset(MemController_4_reset),
    .io_rd_valid(MemController_4_io_rd_valid),
    .io_wr_valid(MemController_4_io_wr_valid),
    .io_rd_data_valid(MemController_4_io_rd_data_valid),
    .io_rd_data_bits(MemController_4_io_rd_data_bits),
    .io_wr_data_valid(MemController_4_io_wr_data_valid),
    .io_wr_data_bits(MemController_4_io_wr_data_bits)
  );
  MemController MemController_5 ( // @[pearray.scala 211:15]
    .clock(MemController_5_clock),
    .reset(MemController_5_reset),
    .io_rd_valid(MemController_5_io_rd_valid),
    .io_wr_valid(MemController_5_io_wr_valid),
    .io_rd_data_valid(MemController_5_io_rd_data_valid),
    .io_rd_data_bits(MemController_5_io_rd_data_bits),
    .io_wr_data_valid(MemController_5_io_wr_data_valid),
    .io_wr_data_bits(MemController_5_io_wr_data_bits)
  );
  MemController MemController_6 ( // @[pearray.scala 211:15]
    .clock(MemController_6_clock),
    .reset(MemController_6_reset),
    .io_rd_valid(MemController_6_io_rd_valid),
    .io_wr_valid(MemController_6_io_wr_valid),
    .io_rd_data_valid(MemController_6_io_rd_data_valid),
    .io_rd_data_bits(MemController_6_io_rd_data_bits),
    .io_wr_data_valid(MemController_6_io_wr_data_valid),
    .io_wr_data_bits(MemController_6_io_wr_data_bits)
  );
  MemController MemController_7 ( // @[pearray.scala 211:15]
    .clock(MemController_7_clock),
    .reset(MemController_7_reset),
    .io_rd_valid(MemController_7_io_rd_valid),
    .io_wr_valid(MemController_7_io_wr_valid),
    .io_rd_data_valid(MemController_7_io_rd_data_valid),
    .io_rd_data_bits(MemController_7_io_rd_data_bits),
    .io_wr_data_valid(MemController_7_io_wr_data_valid),
    .io_wr_data_bits(MemController_7_io_wr_data_bits)
  );
  MemController MemController_8 ( // @[pearray.scala 209:15]
    .clock(MemController_8_clock),
    .reset(MemController_8_reset),
    .io_rd_valid(MemController_8_io_rd_valid),
    .io_wr_valid(MemController_8_io_wr_valid),
    .io_rd_data_valid(MemController_8_io_rd_data_valid),
    .io_rd_data_bits(MemController_8_io_rd_data_bits),
    .io_wr_data_valid(MemController_8_io_wr_data_valid),
    .io_wr_data_bits(MemController_8_io_wr_data_bits)
  );
  MemController MemController_9 ( // @[pearray.scala 209:15]
    .clock(MemController_9_clock),
    .reset(MemController_9_reset),
    .io_rd_valid(MemController_9_io_rd_valid),
    .io_wr_valid(MemController_9_io_wr_valid),
    .io_rd_data_valid(MemController_9_io_rd_data_valid),
    .io_rd_data_bits(MemController_9_io_rd_data_bits),
    .io_wr_data_valid(MemController_9_io_wr_data_valid),
    .io_wr_data_bits(MemController_9_io_wr_data_bits)
  );
  MemController MemController_10 ( // @[pearray.scala 209:15]
    .clock(MemController_10_clock),
    .reset(MemController_10_reset),
    .io_rd_valid(MemController_10_io_rd_valid),
    .io_wr_valid(MemController_10_io_wr_valid),
    .io_rd_data_valid(MemController_10_io_rd_data_valid),
    .io_rd_data_bits(MemController_10_io_rd_data_bits),
    .io_wr_data_valid(MemController_10_io_wr_data_valid),
    .io_wr_data_bits(MemController_10_io_wr_data_bits)
  );
  MemController MemController_11 ( // @[pearray.scala 209:15]
    .clock(MemController_11_clock),
    .reset(MemController_11_reset),
    .io_rd_valid(MemController_11_io_rd_valid),
    .io_wr_valid(MemController_11_io_wr_valid),
    .io_rd_data_valid(MemController_11_io_rd_data_valid),
    .io_rd_data_bits(MemController_11_io_rd_data_bits),
    .io_wr_data_valid(MemController_11_io_wr_data_valid),
    .io_wr_data_bits(MemController_11_io_wr_data_bits)
  );
  MemController MemController_12 ( // @[pearray.scala 209:15]
    .clock(MemController_12_clock),
    .reset(MemController_12_reset),
    .io_rd_valid(MemController_12_io_rd_valid),
    .io_wr_valid(MemController_12_io_wr_valid),
    .io_rd_data_valid(MemController_12_io_rd_data_valid),
    .io_rd_data_bits(MemController_12_io_rd_data_bits),
    .io_wr_data_valid(MemController_12_io_wr_data_valid),
    .io_wr_data_bits(MemController_12_io_wr_data_bits)
  );
  MemController MemController_13 ( // @[pearray.scala 209:15]
    .clock(MemController_13_clock),
    .reset(MemController_13_reset),
    .io_rd_valid(MemController_13_io_rd_valid),
    .io_wr_valid(MemController_13_io_wr_valid),
    .io_rd_data_valid(MemController_13_io_rd_data_valid),
    .io_rd_data_bits(MemController_13_io_rd_data_bits),
    .io_wr_data_valid(MemController_13_io_wr_data_valid),
    .io_wr_data_bits(MemController_13_io_wr_data_bits)
  );
  MemController MemController_14 ( // @[pearray.scala 209:15]
    .clock(MemController_14_clock),
    .reset(MemController_14_reset),
    .io_rd_valid(MemController_14_io_rd_valid),
    .io_wr_valid(MemController_14_io_wr_valid),
    .io_rd_data_valid(MemController_14_io_rd_data_valid),
    .io_rd_data_bits(MemController_14_io_rd_data_bits),
    .io_wr_data_valid(MemController_14_io_wr_data_valid),
    .io_wr_data_bits(MemController_14_io_wr_data_bits)
  );
  MemController MemController_15 ( // @[pearray.scala 209:15]
    .clock(MemController_15_clock),
    .reset(MemController_15_reset),
    .io_rd_valid(MemController_15_io_rd_valid),
    .io_wr_valid(MemController_15_io_wr_valid),
    .io_rd_data_valid(MemController_15_io_rd_data_valid),
    .io_rd_data_bits(MemController_15_io_rd_data_bits),
    .io_wr_data_valid(MemController_15_io_wr_data_valid),
    .io_wr_data_bits(MemController_15_io_wr_data_bits)
  );
  MemController MemController_16 ( // @[pearray.scala 209:15]
    .clock(MemController_16_clock),
    .reset(MemController_16_reset),
    .io_rd_valid(MemController_16_io_rd_valid),
    .io_wr_valid(MemController_16_io_wr_valid),
    .io_rd_data_valid(MemController_16_io_rd_data_valid),
    .io_rd_data_bits(MemController_16_io_rd_data_bits),
    .io_wr_data_valid(MemController_16_io_wr_data_valid),
    .io_wr_data_bits(MemController_16_io_wr_data_bits)
  );
  MemController MemController_17 ( // @[pearray.scala 209:15]
    .clock(MemController_17_clock),
    .reset(MemController_17_reset),
    .io_rd_valid(MemController_17_io_rd_valid),
    .io_wr_valid(MemController_17_io_wr_valid),
    .io_rd_data_valid(MemController_17_io_rd_data_valid),
    .io_rd_data_bits(MemController_17_io_rd_data_bits),
    .io_wr_data_valid(MemController_17_io_wr_data_valid),
    .io_wr_data_bits(MemController_17_io_wr_data_bits)
  );
  MemController MemController_18 ( // @[pearray.scala 209:15]
    .clock(MemController_18_clock),
    .reset(MemController_18_reset),
    .io_rd_valid(MemController_18_io_rd_valid),
    .io_wr_valid(MemController_18_io_wr_valid),
    .io_rd_data_valid(MemController_18_io_rd_data_valid),
    .io_rd_data_bits(MemController_18_io_rd_data_bits),
    .io_wr_data_valid(MemController_18_io_wr_data_valid),
    .io_wr_data_bits(MemController_18_io_wr_data_bits)
  );
  MemController MemController_19 ( // @[pearray.scala 209:15]
    .clock(MemController_19_clock),
    .reset(MemController_19_reset),
    .io_rd_valid(MemController_19_io_rd_valid),
    .io_wr_valid(MemController_19_io_wr_valid),
    .io_rd_data_valid(MemController_19_io_rd_data_valid),
    .io_rd_data_bits(MemController_19_io_rd_data_bits),
    .io_wr_data_valid(MemController_19_io_wr_data_valid),
    .io_wr_data_bits(MemController_19_io_wr_data_bits)
  );
  MemController MemController_20 ( // @[pearray.scala 209:15]
    .clock(MemController_20_clock),
    .reset(MemController_20_reset),
    .io_rd_valid(MemController_20_io_rd_valid),
    .io_wr_valid(MemController_20_io_wr_valid),
    .io_rd_data_valid(MemController_20_io_rd_data_valid),
    .io_rd_data_bits(MemController_20_io_rd_data_bits),
    .io_wr_data_valid(MemController_20_io_wr_data_valid),
    .io_wr_data_bits(MemController_20_io_wr_data_bits)
  );
  MemController MemController_21 ( // @[pearray.scala 209:15]
    .clock(MemController_21_clock),
    .reset(MemController_21_reset),
    .io_rd_valid(MemController_21_io_rd_valid),
    .io_wr_valid(MemController_21_io_wr_valid),
    .io_rd_data_valid(MemController_21_io_rd_data_valid),
    .io_rd_data_bits(MemController_21_io_rd_data_bits),
    .io_wr_data_valid(MemController_21_io_wr_data_valid),
    .io_wr_data_bits(MemController_21_io_wr_data_bits)
  );
  MemController MemController_22 ( // @[pearray.scala 209:15]
    .clock(MemController_22_clock),
    .reset(MemController_22_reset),
    .io_rd_valid(MemController_22_io_rd_valid),
    .io_wr_valid(MemController_22_io_wr_valid),
    .io_rd_data_valid(MemController_22_io_rd_data_valid),
    .io_rd_data_bits(MemController_22_io_rd_data_bits),
    .io_wr_data_valid(MemController_22_io_wr_data_valid),
    .io_wr_data_bits(MemController_22_io_wr_data_bits)
  );
  MemController MemController_23 ( // @[pearray.scala 209:15]
    .clock(MemController_23_clock),
    .reset(MemController_23_reset),
    .io_rd_valid(MemController_23_io_rd_valid),
    .io_wr_valid(MemController_23_io_wr_valid),
    .io_rd_data_valid(MemController_23_io_rd_data_valid),
    .io_rd_data_bits(MemController_23_io_rd_data_bits),
    .io_wr_data_valid(MemController_23_io_wr_data_valid),
    .io_wr_data_bits(MemController_23_io_wr_data_bits)
  );
  assign io_data_0_out_0_valid = MemController_io_rd_data_valid; // @[pearray.scala 256:31]
  assign io_data_0_out_0_bits = MemController_io_rd_data_bits; // @[pearray.scala 256:31]
  assign io_data_0_out_1_valid = MemController_1_io_rd_data_valid; // @[pearray.scala 256:31]
  assign io_data_0_out_1_bits = MemController_1_io_rd_data_bits; // @[pearray.scala 256:31]
  assign io_data_0_out_2_valid = MemController_2_io_rd_data_valid; // @[pearray.scala 256:31]
  assign io_data_0_out_2_bits = MemController_2_io_rd_data_bits; // @[pearray.scala 256:31]
  assign io_data_0_out_3_valid = MemController_3_io_rd_data_valid; // @[pearray.scala 256:31]
  assign io_data_0_out_3_bits = MemController_3_io_rd_data_bits; // @[pearray.scala 256:31]
  assign io_data_0_out_4_valid = MemController_4_io_rd_data_valid; // @[pearray.scala 256:31]
  assign io_data_0_out_4_bits = MemController_4_io_rd_data_bits; // @[pearray.scala 256:31]
  assign io_data_0_out_5_valid = MemController_5_io_rd_data_valid; // @[pearray.scala 256:31]
  assign io_data_0_out_5_bits = MemController_5_io_rd_data_bits; // @[pearray.scala 256:31]
  assign io_data_0_out_6_valid = MemController_6_io_rd_data_valid; // @[pearray.scala 256:31]
  assign io_data_0_out_6_bits = MemController_6_io_rd_data_bits; // @[pearray.scala 256:31]
  assign io_data_0_out_7_valid = MemController_7_io_rd_data_valid; // @[pearray.scala 256:31]
  assign io_data_0_out_7_bits = MemController_7_io_rd_data_bits; // @[pearray.scala 256:31]
  assign MultiDimTime_clock = clock;
  assign MultiDimTime_reset = reset;
  assign MultiDimTime_io_in = io_exec_valid; // @[pearray.scala 149:16]
  assign PE_clock = clock;
  assign PE_reset = reset;
  assign PE_io_data_2_in_valid = PENetwork_16_io_to_pes_0_in_valid; // @[pearray.scala 160:34]
  assign PE_io_data_2_in_bits = PENetwork_16_io_to_pes_0_in_bits; // @[pearray.scala 160:34]
  assign PE_io_data_1_in_valid = PENetwork_8_io_to_pes_0_in_valid; // @[pearray.scala 160:34]
  assign PE_io_data_1_in_bits = PENetwork_8_io_to_pes_0_in_bits; // @[pearray.scala 160:34]
  assign PE_io_data_0_in_valid = 1'h0; // @[pearray.scala 160:34]
  assign PE_io_data_0_in_bits = 16'h0; // @[pearray.scala 160:34]
  assign PE_io_sig_stat2trans = _T_12_3; // @[pearray.scala 184:38]
  assign PE_1_clock = clock;
  assign PE_1_reset = reset;
  assign PE_1_io_data_2_in_valid = PENetwork_17_io_to_pes_0_in_valid; // @[pearray.scala 160:34]
  assign PE_1_io_data_2_in_bits = PENetwork_17_io_to_pes_0_in_bits; // @[pearray.scala 160:34]
  assign PE_1_io_data_1_in_valid = PENetwork_8_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_1_io_data_1_in_bits = PENetwork_8_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_1_io_data_0_in_valid = PENetwork_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_1_io_data_0_in_bits = PENetwork_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_1_io_sig_stat2trans = _T_22_3; // @[pearray.scala 184:38]
  assign PE_2_clock = clock;
  assign PE_2_reset = reset;
  assign PE_2_io_data_2_in_valid = PENetwork_18_io_to_pes_0_in_valid; // @[pearray.scala 160:34]
  assign PE_2_io_data_2_in_bits = PENetwork_18_io_to_pes_0_in_bits; // @[pearray.scala 160:34]
  assign PE_2_io_data_1_in_valid = PENetwork_8_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_2_io_data_1_in_bits = PENetwork_8_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_2_io_data_0_in_valid = PENetwork_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_2_io_data_0_in_bits = PENetwork_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_2_io_sig_stat2trans = _T_32_3; // @[pearray.scala 184:38]
  assign PE_3_clock = clock;
  assign PE_3_reset = reset;
  assign PE_3_io_data_2_in_valid = PENetwork_19_io_to_pes_0_in_valid; // @[pearray.scala 160:34]
  assign PE_3_io_data_2_in_bits = PENetwork_19_io_to_pes_0_in_bits; // @[pearray.scala 160:34]
  assign PE_3_io_data_1_in_valid = PENetwork_8_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_3_io_data_1_in_bits = PENetwork_8_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_3_io_data_0_in_valid = PENetwork_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_3_io_data_0_in_bits = PENetwork_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_3_io_sig_stat2trans = _T_42_3; // @[pearray.scala 184:38]
  assign PE_4_clock = clock;
  assign PE_4_reset = reset;
  assign PE_4_io_data_2_in_valid = PENetwork_20_io_to_pes_0_in_valid; // @[pearray.scala 160:34]
  assign PE_4_io_data_2_in_bits = PENetwork_20_io_to_pes_0_in_bits; // @[pearray.scala 160:34]
  assign PE_4_io_data_1_in_valid = PENetwork_8_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_4_io_data_1_in_bits = PENetwork_8_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_4_io_data_0_in_valid = PENetwork_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_4_io_data_0_in_bits = PENetwork_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_4_io_sig_stat2trans = _T_52_3; // @[pearray.scala 184:38]
  assign PE_5_clock = clock;
  assign PE_5_reset = reset;
  assign PE_5_io_data_2_in_valid = PENetwork_21_io_to_pes_0_in_valid; // @[pearray.scala 160:34]
  assign PE_5_io_data_2_in_bits = PENetwork_21_io_to_pes_0_in_bits; // @[pearray.scala 160:34]
  assign PE_5_io_data_1_in_valid = PENetwork_8_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_5_io_data_1_in_bits = PENetwork_8_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_5_io_data_0_in_valid = PENetwork_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_5_io_data_0_in_bits = PENetwork_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_5_io_sig_stat2trans = _T_62_3; // @[pearray.scala 184:38]
  assign PE_6_clock = clock;
  assign PE_6_reset = reset;
  assign PE_6_io_data_2_in_valid = PENetwork_22_io_to_pes_0_in_valid; // @[pearray.scala 160:34]
  assign PE_6_io_data_2_in_bits = PENetwork_22_io_to_pes_0_in_bits; // @[pearray.scala 160:34]
  assign PE_6_io_data_1_in_valid = PENetwork_8_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_6_io_data_1_in_bits = PENetwork_8_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_6_io_data_0_in_valid = PENetwork_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_6_io_data_0_in_bits = PENetwork_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_6_io_sig_stat2trans = _T_72_3; // @[pearray.scala 184:38]
  assign PE_7_clock = clock;
  assign PE_7_reset = reset;
  assign PE_7_io_data_2_in_valid = PENetwork_23_io_to_pes_0_in_valid; // @[pearray.scala 160:34]
  assign PE_7_io_data_2_in_bits = PENetwork_23_io_to_pes_0_in_bits; // @[pearray.scala 160:34]
  assign PE_7_io_data_1_in_valid = PENetwork_8_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_7_io_data_1_in_bits = PENetwork_8_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_7_io_data_0_in_valid = PENetwork_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_7_io_data_0_in_bits = PENetwork_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_7_io_sig_stat2trans = _T_82_3; // @[pearray.scala 184:38]
  assign PE_8_clock = clock;
  assign PE_8_reset = reset;
  assign PE_8_io_data_2_in_valid = PENetwork_16_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_8_io_data_2_in_bits = PENetwork_16_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_8_io_data_1_in_valid = PENetwork_9_io_to_pes_0_in_valid; // @[pearray.scala 160:34]
  assign PE_8_io_data_1_in_bits = PENetwork_9_io_to_pes_0_in_bits; // @[pearray.scala 160:34]
  assign PE_8_io_data_0_in_valid = 1'h0; // @[pearray.scala 160:34]
  assign PE_8_io_data_0_in_bits = 16'h0; // @[pearray.scala 160:34]
  assign PE_8_io_sig_stat2trans = _T_92_3; // @[pearray.scala 184:38]
  assign PE_9_clock = clock;
  assign PE_9_reset = reset;
  assign PE_9_io_data_2_in_valid = PENetwork_17_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_9_io_data_2_in_bits = PENetwork_17_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_9_io_data_1_in_valid = PENetwork_9_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_9_io_data_1_in_bits = PENetwork_9_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_9_io_data_0_in_valid = PENetwork_1_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_9_io_data_0_in_bits = PENetwork_1_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_9_io_sig_stat2trans = _T_102_3; // @[pearray.scala 184:38]
  assign PE_10_clock = clock;
  assign PE_10_reset = reset;
  assign PE_10_io_data_2_in_valid = PENetwork_18_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_10_io_data_2_in_bits = PENetwork_18_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_10_io_data_1_in_valid = PENetwork_9_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_10_io_data_1_in_bits = PENetwork_9_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_10_io_data_0_in_valid = PENetwork_1_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_10_io_data_0_in_bits = PENetwork_1_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_10_io_sig_stat2trans = _T_112_3; // @[pearray.scala 184:38]
  assign PE_11_clock = clock;
  assign PE_11_reset = reset;
  assign PE_11_io_data_2_in_valid = PENetwork_19_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_11_io_data_2_in_bits = PENetwork_19_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_11_io_data_1_in_valid = PENetwork_9_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_11_io_data_1_in_bits = PENetwork_9_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_11_io_data_0_in_valid = PENetwork_1_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_11_io_data_0_in_bits = PENetwork_1_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_11_io_sig_stat2trans = _T_122_3; // @[pearray.scala 184:38]
  assign PE_12_clock = clock;
  assign PE_12_reset = reset;
  assign PE_12_io_data_2_in_valid = PENetwork_20_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_12_io_data_2_in_bits = PENetwork_20_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_12_io_data_1_in_valid = PENetwork_9_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_12_io_data_1_in_bits = PENetwork_9_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_12_io_data_0_in_valid = PENetwork_1_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_12_io_data_0_in_bits = PENetwork_1_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_12_io_sig_stat2trans = _T_132_3; // @[pearray.scala 184:38]
  assign PE_13_clock = clock;
  assign PE_13_reset = reset;
  assign PE_13_io_data_2_in_valid = PENetwork_21_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_13_io_data_2_in_bits = PENetwork_21_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_13_io_data_1_in_valid = PENetwork_9_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_13_io_data_1_in_bits = PENetwork_9_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_13_io_data_0_in_valid = PENetwork_1_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_13_io_data_0_in_bits = PENetwork_1_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_13_io_sig_stat2trans = _T_142_3; // @[pearray.scala 184:38]
  assign PE_14_clock = clock;
  assign PE_14_reset = reset;
  assign PE_14_io_data_2_in_valid = PENetwork_22_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_14_io_data_2_in_bits = PENetwork_22_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_14_io_data_1_in_valid = PENetwork_9_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_14_io_data_1_in_bits = PENetwork_9_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_14_io_data_0_in_valid = PENetwork_1_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_14_io_data_0_in_bits = PENetwork_1_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_14_io_sig_stat2trans = _T_152_3; // @[pearray.scala 184:38]
  assign PE_15_clock = clock;
  assign PE_15_reset = reset;
  assign PE_15_io_data_2_in_valid = PENetwork_23_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_15_io_data_2_in_bits = PENetwork_23_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_15_io_data_1_in_valid = PENetwork_9_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_15_io_data_1_in_bits = PENetwork_9_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_15_io_data_0_in_valid = PENetwork_1_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_15_io_data_0_in_bits = PENetwork_1_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_15_io_sig_stat2trans = _T_162_3; // @[pearray.scala 184:38]
  assign PE_16_clock = clock;
  assign PE_16_reset = reset;
  assign PE_16_io_data_2_in_valid = PENetwork_16_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_16_io_data_2_in_bits = PENetwork_16_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_16_io_data_1_in_valid = PENetwork_10_io_to_pes_0_in_valid; // @[pearray.scala 160:34]
  assign PE_16_io_data_1_in_bits = PENetwork_10_io_to_pes_0_in_bits; // @[pearray.scala 160:34]
  assign PE_16_io_data_0_in_valid = 1'h0; // @[pearray.scala 160:34]
  assign PE_16_io_data_0_in_bits = 16'h0; // @[pearray.scala 160:34]
  assign PE_16_io_sig_stat2trans = _T_172_3; // @[pearray.scala 184:38]
  assign PE_17_clock = clock;
  assign PE_17_reset = reset;
  assign PE_17_io_data_2_in_valid = PENetwork_17_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_17_io_data_2_in_bits = PENetwork_17_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_17_io_data_1_in_valid = PENetwork_10_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_17_io_data_1_in_bits = PENetwork_10_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_17_io_data_0_in_valid = PENetwork_2_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_17_io_data_0_in_bits = PENetwork_2_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_17_io_sig_stat2trans = _T_182_3; // @[pearray.scala 184:38]
  assign PE_18_clock = clock;
  assign PE_18_reset = reset;
  assign PE_18_io_data_2_in_valid = PENetwork_18_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_18_io_data_2_in_bits = PENetwork_18_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_18_io_data_1_in_valid = PENetwork_10_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_18_io_data_1_in_bits = PENetwork_10_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_18_io_data_0_in_valid = PENetwork_2_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_18_io_data_0_in_bits = PENetwork_2_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_18_io_sig_stat2trans = _T_192_3; // @[pearray.scala 184:38]
  assign PE_19_clock = clock;
  assign PE_19_reset = reset;
  assign PE_19_io_data_2_in_valid = PENetwork_19_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_19_io_data_2_in_bits = PENetwork_19_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_19_io_data_1_in_valid = PENetwork_10_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_19_io_data_1_in_bits = PENetwork_10_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_19_io_data_0_in_valid = PENetwork_2_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_19_io_data_0_in_bits = PENetwork_2_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_19_io_sig_stat2trans = _T_202_3; // @[pearray.scala 184:38]
  assign PE_20_clock = clock;
  assign PE_20_reset = reset;
  assign PE_20_io_data_2_in_valid = PENetwork_20_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_20_io_data_2_in_bits = PENetwork_20_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_20_io_data_1_in_valid = PENetwork_10_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_20_io_data_1_in_bits = PENetwork_10_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_20_io_data_0_in_valid = PENetwork_2_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_20_io_data_0_in_bits = PENetwork_2_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_20_io_sig_stat2trans = _T_212_3; // @[pearray.scala 184:38]
  assign PE_21_clock = clock;
  assign PE_21_reset = reset;
  assign PE_21_io_data_2_in_valid = PENetwork_21_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_21_io_data_2_in_bits = PENetwork_21_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_21_io_data_1_in_valid = PENetwork_10_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_21_io_data_1_in_bits = PENetwork_10_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_21_io_data_0_in_valid = PENetwork_2_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_21_io_data_0_in_bits = PENetwork_2_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_21_io_sig_stat2trans = _T_222_3; // @[pearray.scala 184:38]
  assign PE_22_clock = clock;
  assign PE_22_reset = reset;
  assign PE_22_io_data_2_in_valid = PENetwork_22_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_22_io_data_2_in_bits = PENetwork_22_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_22_io_data_1_in_valid = PENetwork_10_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_22_io_data_1_in_bits = PENetwork_10_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_22_io_data_0_in_valid = PENetwork_2_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_22_io_data_0_in_bits = PENetwork_2_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_22_io_sig_stat2trans = _T_232_3; // @[pearray.scala 184:38]
  assign PE_23_clock = clock;
  assign PE_23_reset = reset;
  assign PE_23_io_data_2_in_valid = PENetwork_23_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_23_io_data_2_in_bits = PENetwork_23_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_23_io_data_1_in_valid = PENetwork_10_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_23_io_data_1_in_bits = PENetwork_10_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_23_io_data_0_in_valid = PENetwork_2_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_23_io_data_0_in_bits = PENetwork_2_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_23_io_sig_stat2trans = _T_242_3; // @[pearray.scala 184:38]
  assign PE_24_clock = clock;
  assign PE_24_reset = reset;
  assign PE_24_io_data_2_in_valid = PENetwork_16_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_24_io_data_2_in_bits = PENetwork_16_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_24_io_data_1_in_valid = PENetwork_11_io_to_pes_0_in_valid; // @[pearray.scala 160:34]
  assign PE_24_io_data_1_in_bits = PENetwork_11_io_to_pes_0_in_bits; // @[pearray.scala 160:34]
  assign PE_24_io_data_0_in_valid = 1'h0; // @[pearray.scala 160:34]
  assign PE_24_io_data_0_in_bits = 16'h0; // @[pearray.scala 160:34]
  assign PE_24_io_sig_stat2trans = _T_252_3; // @[pearray.scala 184:38]
  assign PE_25_clock = clock;
  assign PE_25_reset = reset;
  assign PE_25_io_data_2_in_valid = PENetwork_17_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_25_io_data_2_in_bits = PENetwork_17_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_25_io_data_1_in_valid = PENetwork_11_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_25_io_data_1_in_bits = PENetwork_11_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_25_io_data_0_in_valid = PENetwork_3_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_25_io_data_0_in_bits = PENetwork_3_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_25_io_sig_stat2trans = _T_262_3; // @[pearray.scala 184:38]
  assign PE_26_clock = clock;
  assign PE_26_reset = reset;
  assign PE_26_io_data_2_in_valid = PENetwork_18_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_26_io_data_2_in_bits = PENetwork_18_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_26_io_data_1_in_valid = PENetwork_11_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_26_io_data_1_in_bits = PENetwork_11_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_26_io_data_0_in_valid = PENetwork_3_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_26_io_data_0_in_bits = PENetwork_3_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_26_io_sig_stat2trans = _T_272_3; // @[pearray.scala 184:38]
  assign PE_27_clock = clock;
  assign PE_27_reset = reset;
  assign PE_27_io_data_2_in_valid = PENetwork_19_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_27_io_data_2_in_bits = PENetwork_19_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_27_io_data_1_in_valid = PENetwork_11_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_27_io_data_1_in_bits = PENetwork_11_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_27_io_data_0_in_valid = PENetwork_3_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_27_io_data_0_in_bits = PENetwork_3_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_27_io_sig_stat2trans = _T_282_3; // @[pearray.scala 184:38]
  assign PE_28_clock = clock;
  assign PE_28_reset = reset;
  assign PE_28_io_data_2_in_valid = PENetwork_20_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_28_io_data_2_in_bits = PENetwork_20_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_28_io_data_1_in_valid = PENetwork_11_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_28_io_data_1_in_bits = PENetwork_11_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_28_io_data_0_in_valid = PENetwork_3_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_28_io_data_0_in_bits = PENetwork_3_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_28_io_sig_stat2trans = _T_292_3; // @[pearray.scala 184:38]
  assign PE_29_clock = clock;
  assign PE_29_reset = reset;
  assign PE_29_io_data_2_in_valid = PENetwork_21_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_29_io_data_2_in_bits = PENetwork_21_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_29_io_data_1_in_valid = PENetwork_11_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_29_io_data_1_in_bits = PENetwork_11_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_29_io_data_0_in_valid = PENetwork_3_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_29_io_data_0_in_bits = PENetwork_3_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_29_io_sig_stat2trans = _T_302_3; // @[pearray.scala 184:38]
  assign PE_30_clock = clock;
  assign PE_30_reset = reset;
  assign PE_30_io_data_2_in_valid = PENetwork_22_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_30_io_data_2_in_bits = PENetwork_22_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_30_io_data_1_in_valid = PENetwork_11_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_30_io_data_1_in_bits = PENetwork_11_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_30_io_data_0_in_valid = PENetwork_3_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_30_io_data_0_in_bits = PENetwork_3_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_30_io_sig_stat2trans = _T_312_3; // @[pearray.scala 184:38]
  assign PE_31_clock = clock;
  assign PE_31_reset = reset;
  assign PE_31_io_data_2_in_valid = PENetwork_23_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_31_io_data_2_in_bits = PENetwork_23_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_31_io_data_1_in_valid = PENetwork_11_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_31_io_data_1_in_bits = PENetwork_11_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_31_io_data_0_in_valid = PENetwork_3_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_31_io_data_0_in_bits = PENetwork_3_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_31_io_sig_stat2trans = _T_322_3; // @[pearray.scala 184:38]
  assign PE_32_clock = clock;
  assign PE_32_reset = reset;
  assign PE_32_io_data_2_in_valid = PENetwork_16_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_32_io_data_2_in_bits = PENetwork_16_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_32_io_data_1_in_valid = PENetwork_12_io_to_pes_0_in_valid; // @[pearray.scala 160:34]
  assign PE_32_io_data_1_in_bits = PENetwork_12_io_to_pes_0_in_bits; // @[pearray.scala 160:34]
  assign PE_32_io_data_0_in_valid = 1'h0; // @[pearray.scala 160:34]
  assign PE_32_io_data_0_in_bits = 16'h0; // @[pearray.scala 160:34]
  assign PE_32_io_sig_stat2trans = _T_332_3; // @[pearray.scala 184:38]
  assign PE_33_clock = clock;
  assign PE_33_reset = reset;
  assign PE_33_io_data_2_in_valid = PENetwork_17_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_33_io_data_2_in_bits = PENetwork_17_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_33_io_data_1_in_valid = PENetwork_12_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_33_io_data_1_in_bits = PENetwork_12_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_33_io_data_0_in_valid = PENetwork_4_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_33_io_data_0_in_bits = PENetwork_4_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_33_io_sig_stat2trans = _T_342_3; // @[pearray.scala 184:38]
  assign PE_34_clock = clock;
  assign PE_34_reset = reset;
  assign PE_34_io_data_2_in_valid = PENetwork_18_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_34_io_data_2_in_bits = PENetwork_18_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_34_io_data_1_in_valid = PENetwork_12_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_34_io_data_1_in_bits = PENetwork_12_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_34_io_data_0_in_valid = PENetwork_4_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_34_io_data_0_in_bits = PENetwork_4_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_34_io_sig_stat2trans = _T_352_3; // @[pearray.scala 184:38]
  assign PE_35_clock = clock;
  assign PE_35_reset = reset;
  assign PE_35_io_data_2_in_valid = PENetwork_19_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_35_io_data_2_in_bits = PENetwork_19_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_35_io_data_1_in_valid = PENetwork_12_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_35_io_data_1_in_bits = PENetwork_12_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_35_io_data_0_in_valid = PENetwork_4_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_35_io_data_0_in_bits = PENetwork_4_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_35_io_sig_stat2trans = _T_362_3; // @[pearray.scala 184:38]
  assign PE_36_clock = clock;
  assign PE_36_reset = reset;
  assign PE_36_io_data_2_in_valid = PENetwork_20_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_36_io_data_2_in_bits = PENetwork_20_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_36_io_data_1_in_valid = PENetwork_12_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_36_io_data_1_in_bits = PENetwork_12_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_36_io_data_0_in_valid = PENetwork_4_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_36_io_data_0_in_bits = PENetwork_4_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_36_io_sig_stat2trans = _T_372_3; // @[pearray.scala 184:38]
  assign PE_37_clock = clock;
  assign PE_37_reset = reset;
  assign PE_37_io_data_2_in_valid = PENetwork_21_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_37_io_data_2_in_bits = PENetwork_21_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_37_io_data_1_in_valid = PENetwork_12_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_37_io_data_1_in_bits = PENetwork_12_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_37_io_data_0_in_valid = PENetwork_4_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_37_io_data_0_in_bits = PENetwork_4_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_37_io_sig_stat2trans = _T_382_3; // @[pearray.scala 184:38]
  assign PE_38_clock = clock;
  assign PE_38_reset = reset;
  assign PE_38_io_data_2_in_valid = PENetwork_22_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_38_io_data_2_in_bits = PENetwork_22_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_38_io_data_1_in_valid = PENetwork_12_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_38_io_data_1_in_bits = PENetwork_12_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_38_io_data_0_in_valid = PENetwork_4_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_38_io_data_0_in_bits = PENetwork_4_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_38_io_sig_stat2trans = _T_392_3; // @[pearray.scala 184:38]
  assign PE_39_clock = clock;
  assign PE_39_reset = reset;
  assign PE_39_io_data_2_in_valid = PENetwork_23_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_39_io_data_2_in_bits = PENetwork_23_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_39_io_data_1_in_valid = PENetwork_12_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_39_io_data_1_in_bits = PENetwork_12_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_39_io_data_0_in_valid = PENetwork_4_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_39_io_data_0_in_bits = PENetwork_4_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_39_io_sig_stat2trans = _T_402_3; // @[pearray.scala 184:38]
  assign PE_40_clock = clock;
  assign PE_40_reset = reset;
  assign PE_40_io_data_2_in_valid = PENetwork_16_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_40_io_data_2_in_bits = PENetwork_16_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_40_io_data_1_in_valid = PENetwork_13_io_to_pes_0_in_valid; // @[pearray.scala 160:34]
  assign PE_40_io_data_1_in_bits = PENetwork_13_io_to_pes_0_in_bits; // @[pearray.scala 160:34]
  assign PE_40_io_data_0_in_valid = 1'h0; // @[pearray.scala 160:34]
  assign PE_40_io_data_0_in_bits = 16'h0; // @[pearray.scala 160:34]
  assign PE_40_io_sig_stat2trans = _T_412_3; // @[pearray.scala 184:38]
  assign PE_41_clock = clock;
  assign PE_41_reset = reset;
  assign PE_41_io_data_2_in_valid = PENetwork_17_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_41_io_data_2_in_bits = PENetwork_17_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_41_io_data_1_in_valid = PENetwork_13_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_41_io_data_1_in_bits = PENetwork_13_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_41_io_data_0_in_valid = PENetwork_5_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_41_io_data_0_in_bits = PENetwork_5_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_41_io_sig_stat2trans = _T_422_3; // @[pearray.scala 184:38]
  assign PE_42_clock = clock;
  assign PE_42_reset = reset;
  assign PE_42_io_data_2_in_valid = PENetwork_18_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_42_io_data_2_in_bits = PENetwork_18_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_42_io_data_1_in_valid = PENetwork_13_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_42_io_data_1_in_bits = PENetwork_13_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_42_io_data_0_in_valid = PENetwork_5_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_42_io_data_0_in_bits = PENetwork_5_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_42_io_sig_stat2trans = _T_432_3; // @[pearray.scala 184:38]
  assign PE_43_clock = clock;
  assign PE_43_reset = reset;
  assign PE_43_io_data_2_in_valid = PENetwork_19_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_43_io_data_2_in_bits = PENetwork_19_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_43_io_data_1_in_valid = PENetwork_13_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_43_io_data_1_in_bits = PENetwork_13_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_43_io_data_0_in_valid = PENetwork_5_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_43_io_data_0_in_bits = PENetwork_5_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_43_io_sig_stat2trans = _T_442_3; // @[pearray.scala 184:38]
  assign PE_44_clock = clock;
  assign PE_44_reset = reset;
  assign PE_44_io_data_2_in_valid = PENetwork_20_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_44_io_data_2_in_bits = PENetwork_20_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_44_io_data_1_in_valid = PENetwork_13_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_44_io_data_1_in_bits = PENetwork_13_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_44_io_data_0_in_valid = PENetwork_5_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_44_io_data_0_in_bits = PENetwork_5_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_44_io_sig_stat2trans = _T_452_3; // @[pearray.scala 184:38]
  assign PE_45_clock = clock;
  assign PE_45_reset = reset;
  assign PE_45_io_data_2_in_valid = PENetwork_21_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_45_io_data_2_in_bits = PENetwork_21_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_45_io_data_1_in_valid = PENetwork_13_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_45_io_data_1_in_bits = PENetwork_13_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_45_io_data_0_in_valid = PENetwork_5_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_45_io_data_0_in_bits = PENetwork_5_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_45_io_sig_stat2trans = _T_462_3; // @[pearray.scala 184:38]
  assign PE_46_clock = clock;
  assign PE_46_reset = reset;
  assign PE_46_io_data_2_in_valid = PENetwork_22_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_46_io_data_2_in_bits = PENetwork_22_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_46_io_data_1_in_valid = PENetwork_13_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_46_io_data_1_in_bits = PENetwork_13_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_46_io_data_0_in_valid = PENetwork_5_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_46_io_data_0_in_bits = PENetwork_5_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_46_io_sig_stat2trans = _T_472_3; // @[pearray.scala 184:38]
  assign PE_47_clock = clock;
  assign PE_47_reset = reset;
  assign PE_47_io_data_2_in_valid = PENetwork_23_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_47_io_data_2_in_bits = PENetwork_23_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_47_io_data_1_in_valid = PENetwork_13_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_47_io_data_1_in_bits = PENetwork_13_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_47_io_data_0_in_valid = PENetwork_5_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_47_io_data_0_in_bits = PENetwork_5_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_47_io_sig_stat2trans = _T_482_3; // @[pearray.scala 184:38]
  assign PE_48_clock = clock;
  assign PE_48_reset = reset;
  assign PE_48_io_data_2_in_valid = PENetwork_16_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_48_io_data_2_in_bits = PENetwork_16_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_48_io_data_1_in_valid = PENetwork_14_io_to_pes_0_in_valid; // @[pearray.scala 160:34]
  assign PE_48_io_data_1_in_bits = PENetwork_14_io_to_pes_0_in_bits; // @[pearray.scala 160:34]
  assign PE_48_io_data_0_in_valid = 1'h0; // @[pearray.scala 160:34]
  assign PE_48_io_data_0_in_bits = 16'h0; // @[pearray.scala 160:34]
  assign PE_48_io_sig_stat2trans = _T_492_3; // @[pearray.scala 184:38]
  assign PE_49_clock = clock;
  assign PE_49_reset = reset;
  assign PE_49_io_data_2_in_valid = PENetwork_17_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_49_io_data_2_in_bits = PENetwork_17_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_49_io_data_1_in_valid = PENetwork_14_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_49_io_data_1_in_bits = PENetwork_14_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_49_io_data_0_in_valid = PENetwork_6_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_49_io_data_0_in_bits = PENetwork_6_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_49_io_sig_stat2trans = _T_502_3; // @[pearray.scala 184:38]
  assign PE_50_clock = clock;
  assign PE_50_reset = reset;
  assign PE_50_io_data_2_in_valid = PENetwork_18_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_50_io_data_2_in_bits = PENetwork_18_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_50_io_data_1_in_valid = PENetwork_14_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_50_io_data_1_in_bits = PENetwork_14_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_50_io_data_0_in_valid = PENetwork_6_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_50_io_data_0_in_bits = PENetwork_6_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_50_io_sig_stat2trans = _T_512_3; // @[pearray.scala 184:38]
  assign PE_51_clock = clock;
  assign PE_51_reset = reset;
  assign PE_51_io_data_2_in_valid = PENetwork_19_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_51_io_data_2_in_bits = PENetwork_19_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_51_io_data_1_in_valid = PENetwork_14_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_51_io_data_1_in_bits = PENetwork_14_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_51_io_data_0_in_valid = PENetwork_6_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_51_io_data_0_in_bits = PENetwork_6_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_51_io_sig_stat2trans = _T_522_3; // @[pearray.scala 184:38]
  assign PE_52_clock = clock;
  assign PE_52_reset = reset;
  assign PE_52_io_data_2_in_valid = PENetwork_20_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_52_io_data_2_in_bits = PENetwork_20_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_52_io_data_1_in_valid = PENetwork_14_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_52_io_data_1_in_bits = PENetwork_14_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_52_io_data_0_in_valid = PENetwork_6_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_52_io_data_0_in_bits = PENetwork_6_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_52_io_sig_stat2trans = _T_532_3; // @[pearray.scala 184:38]
  assign PE_53_clock = clock;
  assign PE_53_reset = reset;
  assign PE_53_io_data_2_in_valid = PENetwork_21_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_53_io_data_2_in_bits = PENetwork_21_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_53_io_data_1_in_valid = PENetwork_14_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_53_io_data_1_in_bits = PENetwork_14_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_53_io_data_0_in_valid = PENetwork_6_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_53_io_data_0_in_bits = PENetwork_6_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_53_io_sig_stat2trans = _T_542_3; // @[pearray.scala 184:38]
  assign PE_54_clock = clock;
  assign PE_54_reset = reset;
  assign PE_54_io_data_2_in_valid = PENetwork_22_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_54_io_data_2_in_bits = PENetwork_22_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_54_io_data_1_in_valid = PENetwork_14_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_54_io_data_1_in_bits = PENetwork_14_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_54_io_data_0_in_valid = PENetwork_6_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_54_io_data_0_in_bits = PENetwork_6_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_54_io_sig_stat2trans = _T_552_3; // @[pearray.scala 184:38]
  assign PE_55_clock = clock;
  assign PE_55_reset = reset;
  assign PE_55_io_data_2_in_valid = PENetwork_23_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_55_io_data_2_in_bits = PENetwork_23_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_55_io_data_1_in_valid = PENetwork_14_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_55_io_data_1_in_bits = PENetwork_14_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_55_io_data_0_in_valid = PENetwork_6_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_55_io_data_0_in_bits = PENetwork_6_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_55_io_sig_stat2trans = _T_562_3; // @[pearray.scala 184:38]
  assign PE_56_clock = clock;
  assign PE_56_reset = reset;
  assign PE_56_io_data_2_in_valid = PENetwork_16_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_56_io_data_2_in_bits = PENetwork_16_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_56_io_data_1_in_valid = PENetwork_15_io_to_pes_0_in_valid; // @[pearray.scala 160:34]
  assign PE_56_io_data_1_in_bits = PENetwork_15_io_to_pes_0_in_bits; // @[pearray.scala 160:34]
  assign PE_56_io_data_0_in_valid = 1'h0; // @[pearray.scala 160:34]
  assign PE_56_io_data_0_in_bits = 16'h0; // @[pearray.scala 160:34]
  assign PE_56_io_sig_stat2trans = _T_572_3; // @[pearray.scala 184:38]
  assign PE_57_clock = clock;
  assign PE_57_reset = reset;
  assign PE_57_io_data_2_in_valid = PENetwork_17_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_57_io_data_2_in_bits = PENetwork_17_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_57_io_data_1_in_valid = PENetwork_15_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_57_io_data_1_in_bits = PENetwork_15_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_57_io_data_0_in_valid = PENetwork_7_io_to_pes_1_in_valid; // @[pearray.scala 160:34]
  assign PE_57_io_data_0_in_bits = PENetwork_7_io_to_pes_1_in_bits; // @[pearray.scala 160:34]
  assign PE_57_io_sig_stat2trans = _T_582_3; // @[pearray.scala 184:38]
  assign PE_58_clock = clock;
  assign PE_58_reset = reset;
  assign PE_58_io_data_2_in_valid = PENetwork_18_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_58_io_data_2_in_bits = PENetwork_18_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_58_io_data_1_in_valid = PENetwork_15_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_58_io_data_1_in_bits = PENetwork_15_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_58_io_data_0_in_valid = PENetwork_7_io_to_pes_2_in_valid; // @[pearray.scala 160:34]
  assign PE_58_io_data_0_in_bits = PENetwork_7_io_to_pes_2_in_bits; // @[pearray.scala 160:34]
  assign PE_58_io_sig_stat2trans = _T_592_3; // @[pearray.scala 184:38]
  assign PE_59_clock = clock;
  assign PE_59_reset = reset;
  assign PE_59_io_data_2_in_valid = PENetwork_19_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_59_io_data_2_in_bits = PENetwork_19_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_59_io_data_1_in_valid = PENetwork_15_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_59_io_data_1_in_bits = PENetwork_15_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_59_io_data_0_in_valid = PENetwork_7_io_to_pes_3_in_valid; // @[pearray.scala 160:34]
  assign PE_59_io_data_0_in_bits = PENetwork_7_io_to_pes_3_in_bits; // @[pearray.scala 160:34]
  assign PE_59_io_sig_stat2trans = _T_602_3; // @[pearray.scala 184:38]
  assign PE_60_clock = clock;
  assign PE_60_reset = reset;
  assign PE_60_io_data_2_in_valid = PENetwork_20_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_60_io_data_2_in_bits = PENetwork_20_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_60_io_data_1_in_valid = PENetwork_15_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_60_io_data_1_in_bits = PENetwork_15_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_60_io_data_0_in_valid = PENetwork_7_io_to_pes_4_in_valid; // @[pearray.scala 160:34]
  assign PE_60_io_data_0_in_bits = PENetwork_7_io_to_pes_4_in_bits; // @[pearray.scala 160:34]
  assign PE_60_io_sig_stat2trans = _T_612_3; // @[pearray.scala 184:38]
  assign PE_61_clock = clock;
  assign PE_61_reset = reset;
  assign PE_61_io_data_2_in_valid = PENetwork_21_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_61_io_data_2_in_bits = PENetwork_21_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_61_io_data_1_in_valid = PENetwork_15_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_61_io_data_1_in_bits = PENetwork_15_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_61_io_data_0_in_valid = PENetwork_7_io_to_pes_5_in_valid; // @[pearray.scala 160:34]
  assign PE_61_io_data_0_in_bits = PENetwork_7_io_to_pes_5_in_bits; // @[pearray.scala 160:34]
  assign PE_61_io_sig_stat2trans = _T_622_3; // @[pearray.scala 184:38]
  assign PE_62_clock = clock;
  assign PE_62_reset = reset;
  assign PE_62_io_data_2_in_valid = PENetwork_22_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_62_io_data_2_in_bits = PENetwork_22_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_62_io_data_1_in_valid = PENetwork_15_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_62_io_data_1_in_bits = PENetwork_15_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_62_io_data_0_in_valid = PENetwork_7_io_to_pes_6_in_valid; // @[pearray.scala 160:34]
  assign PE_62_io_data_0_in_bits = PENetwork_7_io_to_pes_6_in_bits; // @[pearray.scala 160:34]
  assign PE_62_io_sig_stat2trans = _T_632_3; // @[pearray.scala 184:38]
  assign PE_63_clock = clock;
  assign PE_63_reset = reset;
  assign PE_63_io_data_2_in_valid = PENetwork_23_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_63_io_data_2_in_bits = PENetwork_23_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_63_io_data_1_in_valid = PENetwork_15_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_63_io_data_1_in_bits = PENetwork_15_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_63_io_data_0_in_valid = PENetwork_7_io_to_pes_7_in_valid; // @[pearray.scala 160:34]
  assign PE_63_io_data_0_in_bits = PENetwork_7_io_to_pes_7_in_bits; // @[pearray.scala 160:34]
  assign PE_63_io_sig_stat2trans = _T_642_3; // @[pearray.scala 184:38]
  assign PENetwork_io_to_pes_0_out_valid = PE_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_io_to_pes_0_out_bits = PE_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_io_to_pes_1_out_valid = PE_1_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_io_to_pes_1_out_bits = PE_1_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_io_to_pes_2_out_valid = PE_2_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_io_to_pes_2_out_bits = PE_2_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_io_to_pes_3_out_valid = PE_3_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_io_to_pes_3_out_bits = PE_3_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_io_to_pes_4_out_valid = PE_4_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_io_to_pes_4_out_bits = PE_4_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_io_to_pes_5_out_valid = PE_5_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_io_to_pes_5_out_bits = PE_5_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_io_to_pes_6_out_valid = PE_6_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_io_to_pes_6_out_bits = PE_6_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_io_to_pes_7_out_valid = PE_7_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_io_to_pes_7_out_bits = PE_7_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_1_io_to_pes_0_out_valid = PE_8_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_1_io_to_pes_0_out_bits = PE_8_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_1_io_to_pes_1_out_valid = PE_9_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_1_io_to_pes_1_out_bits = PE_9_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_1_io_to_pes_2_out_valid = PE_10_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_1_io_to_pes_2_out_bits = PE_10_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_1_io_to_pes_3_out_valid = PE_11_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_1_io_to_pes_3_out_bits = PE_11_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_1_io_to_pes_4_out_valid = PE_12_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_1_io_to_pes_4_out_bits = PE_12_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_1_io_to_pes_5_out_valid = PE_13_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_1_io_to_pes_5_out_bits = PE_13_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_1_io_to_pes_6_out_valid = PE_14_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_1_io_to_pes_6_out_bits = PE_14_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_1_io_to_pes_7_out_valid = PE_15_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_1_io_to_pes_7_out_bits = PE_15_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_2_io_to_pes_0_out_valid = PE_16_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_2_io_to_pes_0_out_bits = PE_16_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_2_io_to_pes_1_out_valid = PE_17_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_2_io_to_pes_1_out_bits = PE_17_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_2_io_to_pes_2_out_valid = PE_18_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_2_io_to_pes_2_out_bits = PE_18_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_2_io_to_pes_3_out_valid = PE_19_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_2_io_to_pes_3_out_bits = PE_19_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_2_io_to_pes_4_out_valid = PE_20_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_2_io_to_pes_4_out_bits = PE_20_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_2_io_to_pes_5_out_valid = PE_21_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_2_io_to_pes_5_out_bits = PE_21_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_2_io_to_pes_6_out_valid = PE_22_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_2_io_to_pes_6_out_bits = PE_22_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_2_io_to_pes_7_out_valid = PE_23_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_2_io_to_pes_7_out_bits = PE_23_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_3_io_to_pes_0_out_valid = PE_24_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_3_io_to_pes_0_out_bits = PE_24_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_3_io_to_pes_1_out_valid = PE_25_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_3_io_to_pes_1_out_bits = PE_25_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_3_io_to_pes_2_out_valid = PE_26_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_3_io_to_pes_2_out_bits = PE_26_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_3_io_to_pes_3_out_valid = PE_27_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_3_io_to_pes_3_out_bits = PE_27_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_3_io_to_pes_4_out_valid = PE_28_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_3_io_to_pes_4_out_bits = PE_28_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_3_io_to_pes_5_out_valid = PE_29_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_3_io_to_pes_5_out_bits = PE_29_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_3_io_to_pes_6_out_valid = PE_30_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_3_io_to_pes_6_out_bits = PE_30_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_3_io_to_pes_7_out_valid = PE_31_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_3_io_to_pes_7_out_bits = PE_31_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_4_io_to_pes_0_out_valid = PE_32_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_4_io_to_pes_0_out_bits = PE_32_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_4_io_to_pes_1_out_valid = PE_33_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_4_io_to_pes_1_out_bits = PE_33_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_4_io_to_pes_2_out_valid = PE_34_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_4_io_to_pes_2_out_bits = PE_34_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_4_io_to_pes_3_out_valid = PE_35_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_4_io_to_pes_3_out_bits = PE_35_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_4_io_to_pes_4_out_valid = PE_36_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_4_io_to_pes_4_out_bits = PE_36_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_4_io_to_pes_5_out_valid = PE_37_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_4_io_to_pes_5_out_bits = PE_37_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_4_io_to_pes_6_out_valid = PE_38_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_4_io_to_pes_6_out_bits = PE_38_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_4_io_to_pes_7_out_valid = PE_39_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_4_io_to_pes_7_out_bits = PE_39_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_5_io_to_pes_0_out_valid = PE_40_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_5_io_to_pes_0_out_bits = PE_40_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_5_io_to_pes_1_out_valid = PE_41_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_5_io_to_pes_1_out_bits = PE_41_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_5_io_to_pes_2_out_valid = PE_42_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_5_io_to_pes_2_out_bits = PE_42_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_5_io_to_pes_3_out_valid = PE_43_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_5_io_to_pes_3_out_bits = PE_43_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_5_io_to_pes_4_out_valid = PE_44_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_5_io_to_pes_4_out_bits = PE_44_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_5_io_to_pes_5_out_valid = PE_45_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_5_io_to_pes_5_out_bits = PE_45_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_5_io_to_pes_6_out_valid = PE_46_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_5_io_to_pes_6_out_bits = PE_46_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_5_io_to_pes_7_out_valid = PE_47_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_5_io_to_pes_7_out_bits = PE_47_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_6_io_to_pes_0_out_valid = PE_48_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_6_io_to_pes_0_out_bits = PE_48_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_6_io_to_pes_1_out_valid = PE_49_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_6_io_to_pes_1_out_bits = PE_49_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_6_io_to_pes_2_out_valid = PE_50_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_6_io_to_pes_2_out_bits = PE_50_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_6_io_to_pes_3_out_valid = PE_51_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_6_io_to_pes_3_out_bits = PE_51_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_6_io_to_pes_4_out_valid = PE_52_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_6_io_to_pes_4_out_bits = PE_52_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_6_io_to_pes_5_out_valid = PE_53_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_6_io_to_pes_5_out_bits = PE_53_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_6_io_to_pes_6_out_valid = PE_54_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_6_io_to_pes_6_out_bits = PE_54_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_6_io_to_pes_7_out_valid = PE_55_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_6_io_to_pes_7_out_bits = PE_55_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_7_io_to_pes_0_out_valid = PE_56_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_7_io_to_pes_0_out_bits = PE_56_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_7_io_to_pes_1_out_valid = PE_57_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_7_io_to_pes_1_out_bits = PE_57_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_7_io_to_pes_2_out_valid = PE_58_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_7_io_to_pes_2_out_bits = PE_58_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_7_io_to_pes_3_out_valid = PE_59_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_7_io_to_pes_3_out_bits = PE_59_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_7_io_to_pes_4_out_valid = PE_60_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_7_io_to_pes_4_out_bits = PE_60_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_7_io_to_pes_5_out_valid = PE_61_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_7_io_to_pes_5_out_bits = PE_61_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_7_io_to_pes_6_out_valid = PE_62_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_7_io_to_pes_6_out_bits = PE_62_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_7_io_to_pes_7_out_valid = PE_63_io_data_0_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_7_io_to_pes_7_out_bits = PE_63_io_data_0_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_8_io_to_pes_0_out_valid = PE_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_8_io_to_pes_0_out_bits = PE_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_8_io_to_pes_1_out_valid = PE_1_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_8_io_to_pes_1_out_bits = PE_1_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_8_io_to_pes_2_out_valid = PE_2_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_8_io_to_pes_2_out_bits = PE_2_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_8_io_to_pes_3_out_valid = PE_3_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_8_io_to_pes_3_out_bits = PE_3_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_8_io_to_pes_4_out_valid = PE_4_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_8_io_to_pes_4_out_bits = PE_4_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_8_io_to_pes_5_out_valid = PE_5_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_8_io_to_pes_5_out_bits = PE_5_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_8_io_to_pes_6_out_valid = PE_6_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_8_io_to_pes_6_out_bits = PE_6_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_8_io_to_mem_valid = MemController_8_io_rd_data_valid; // @[pearray.scala 251:29]
  assign PENetwork_8_io_to_mem_bits = MemController_8_io_rd_data_bits; // @[pearray.scala 251:29]
  assign PENetwork_9_io_to_pes_0_out_valid = PE_8_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_9_io_to_pes_0_out_bits = PE_8_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_9_io_to_pes_1_out_valid = PE_9_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_9_io_to_pes_1_out_bits = PE_9_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_9_io_to_pes_2_out_valid = PE_10_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_9_io_to_pes_2_out_bits = PE_10_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_9_io_to_pes_3_out_valid = PE_11_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_9_io_to_pes_3_out_bits = PE_11_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_9_io_to_pes_4_out_valid = PE_12_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_9_io_to_pes_4_out_bits = PE_12_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_9_io_to_pes_5_out_valid = PE_13_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_9_io_to_pes_5_out_bits = PE_13_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_9_io_to_pes_6_out_valid = PE_14_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_9_io_to_pes_6_out_bits = PE_14_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_9_io_to_mem_valid = MemController_9_io_rd_data_valid; // @[pearray.scala 251:29]
  assign PENetwork_9_io_to_mem_bits = MemController_9_io_rd_data_bits; // @[pearray.scala 251:29]
  assign PENetwork_10_io_to_pes_0_out_valid = PE_16_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_10_io_to_pes_0_out_bits = PE_16_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_10_io_to_pes_1_out_valid = PE_17_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_10_io_to_pes_1_out_bits = PE_17_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_10_io_to_pes_2_out_valid = PE_18_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_10_io_to_pes_2_out_bits = PE_18_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_10_io_to_pes_3_out_valid = PE_19_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_10_io_to_pes_3_out_bits = PE_19_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_10_io_to_pes_4_out_valid = PE_20_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_10_io_to_pes_4_out_bits = PE_20_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_10_io_to_pes_5_out_valid = PE_21_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_10_io_to_pes_5_out_bits = PE_21_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_10_io_to_pes_6_out_valid = PE_22_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_10_io_to_pes_6_out_bits = PE_22_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_10_io_to_mem_valid = MemController_10_io_rd_data_valid; // @[pearray.scala 251:29]
  assign PENetwork_10_io_to_mem_bits = MemController_10_io_rd_data_bits; // @[pearray.scala 251:29]
  assign PENetwork_11_io_to_pes_0_out_valid = PE_24_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_11_io_to_pes_0_out_bits = PE_24_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_11_io_to_pes_1_out_valid = PE_25_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_11_io_to_pes_1_out_bits = PE_25_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_11_io_to_pes_2_out_valid = PE_26_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_11_io_to_pes_2_out_bits = PE_26_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_11_io_to_pes_3_out_valid = PE_27_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_11_io_to_pes_3_out_bits = PE_27_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_11_io_to_pes_4_out_valid = PE_28_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_11_io_to_pes_4_out_bits = PE_28_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_11_io_to_pes_5_out_valid = PE_29_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_11_io_to_pes_5_out_bits = PE_29_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_11_io_to_pes_6_out_valid = PE_30_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_11_io_to_pes_6_out_bits = PE_30_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_11_io_to_mem_valid = MemController_11_io_rd_data_valid; // @[pearray.scala 251:29]
  assign PENetwork_11_io_to_mem_bits = MemController_11_io_rd_data_bits; // @[pearray.scala 251:29]
  assign PENetwork_12_io_to_pes_0_out_valid = PE_32_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_12_io_to_pes_0_out_bits = PE_32_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_12_io_to_pes_1_out_valid = PE_33_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_12_io_to_pes_1_out_bits = PE_33_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_12_io_to_pes_2_out_valid = PE_34_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_12_io_to_pes_2_out_bits = PE_34_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_12_io_to_pes_3_out_valid = PE_35_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_12_io_to_pes_3_out_bits = PE_35_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_12_io_to_pes_4_out_valid = PE_36_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_12_io_to_pes_4_out_bits = PE_36_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_12_io_to_pes_5_out_valid = PE_37_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_12_io_to_pes_5_out_bits = PE_37_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_12_io_to_pes_6_out_valid = PE_38_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_12_io_to_pes_6_out_bits = PE_38_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_12_io_to_mem_valid = MemController_12_io_rd_data_valid; // @[pearray.scala 251:29]
  assign PENetwork_12_io_to_mem_bits = MemController_12_io_rd_data_bits; // @[pearray.scala 251:29]
  assign PENetwork_13_io_to_pes_0_out_valid = PE_40_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_13_io_to_pes_0_out_bits = PE_40_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_13_io_to_pes_1_out_valid = PE_41_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_13_io_to_pes_1_out_bits = PE_41_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_13_io_to_pes_2_out_valid = PE_42_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_13_io_to_pes_2_out_bits = PE_42_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_13_io_to_pes_3_out_valid = PE_43_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_13_io_to_pes_3_out_bits = PE_43_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_13_io_to_pes_4_out_valid = PE_44_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_13_io_to_pes_4_out_bits = PE_44_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_13_io_to_pes_5_out_valid = PE_45_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_13_io_to_pes_5_out_bits = PE_45_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_13_io_to_pes_6_out_valid = PE_46_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_13_io_to_pes_6_out_bits = PE_46_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_13_io_to_mem_valid = MemController_13_io_rd_data_valid; // @[pearray.scala 251:29]
  assign PENetwork_13_io_to_mem_bits = MemController_13_io_rd_data_bits; // @[pearray.scala 251:29]
  assign PENetwork_14_io_to_pes_0_out_valid = PE_48_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_14_io_to_pes_0_out_bits = PE_48_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_14_io_to_pes_1_out_valid = PE_49_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_14_io_to_pes_1_out_bits = PE_49_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_14_io_to_pes_2_out_valid = PE_50_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_14_io_to_pes_2_out_bits = PE_50_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_14_io_to_pes_3_out_valid = PE_51_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_14_io_to_pes_3_out_bits = PE_51_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_14_io_to_pes_4_out_valid = PE_52_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_14_io_to_pes_4_out_bits = PE_52_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_14_io_to_pes_5_out_valid = PE_53_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_14_io_to_pes_5_out_bits = PE_53_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_14_io_to_pes_6_out_valid = PE_54_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_14_io_to_pes_6_out_bits = PE_54_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_14_io_to_mem_valid = MemController_14_io_rd_data_valid; // @[pearray.scala 251:29]
  assign PENetwork_14_io_to_mem_bits = MemController_14_io_rd_data_bits; // @[pearray.scala 251:29]
  assign PENetwork_15_io_to_pes_0_out_valid = PE_56_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_15_io_to_pes_0_out_bits = PE_56_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_15_io_to_pes_1_out_valid = PE_57_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_15_io_to_pes_1_out_bits = PE_57_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_15_io_to_pes_2_out_valid = PE_58_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_15_io_to_pes_2_out_bits = PE_58_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_15_io_to_pes_3_out_valid = PE_59_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_15_io_to_pes_3_out_bits = PE_59_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_15_io_to_pes_4_out_valid = PE_60_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_15_io_to_pes_4_out_bits = PE_60_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_15_io_to_pes_5_out_valid = PE_61_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_15_io_to_pes_5_out_bits = PE_61_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_15_io_to_pes_6_out_valid = PE_62_io_data_1_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_15_io_to_pes_6_out_bits = PE_62_io_data_1_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_15_io_to_mem_valid = MemController_15_io_rd_data_valid; // @[pearray.scala 251:29]
  assign PENetwork_15_io_to_mem_bits = MemController_15_io_rd_data_bits; // @[pearray.scala 251:29]
  assign PENetwork_16_io_to_pes_0_out_valid = PE_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_16_io_to_pes_0_out_bits = PE_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_16_io_to_pes_1_out_valid = PE_8_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_16_io_to_pes_1_out_bits = PE_8_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_16_io_to_pes_2_out_valid = PE_16_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_16_io_to_pes_2_out_bits = PE_16_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_16_io_to_pes_3_out_valid = PE_24_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_16_io_to_pes_3_out_bits = PE_24_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_16_io_to_pes_4_out_valid = PE_32_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_16_io_to_pes_4_out_bits = PE_32_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_16_io_to_pes_5_out_valid = PE_40_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_16_io_to_pes_5_out_bits = PE_40_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_16_io_to_pes_6_out_valid = PE_48_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_16_io_to_pes_6_out_bits = PE_48_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_16_io_to_mem_valid = MemController_16_io_rd_data_valid; // @[pearray.scala 251:29]
  assign PENetwork_16_io_to_mem_bits = MemController_16_io_rd_data_bits; // @[pearray.scala 251:29]
  assign PENetwork_17_io_to_pes_0_out_valid = PE_1_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_17_io_to_pes_0_out_bits = PE_1_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_17_io_to_pes_1_out_valid = PE_9_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_17_io_to_pes_1_out_bits = PE_9_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_17_io_to_pes_2_out_valid = PE_17_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_17_io_to_pes_2_out_bits = PE_17_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_17_io_to_pes_3_out_valid = PE_25_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_17_io_to_pes_3_out_bits = PE_25_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_17_io_to_pes_4_out_valid = PE_33_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_17_io_to_pes_4_out_bits = PE_33_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_17_io_to_pes_5_out_valid = PE_41_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_17_io_to_pes_5_out_bits = PE_41_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_17_io_to_pes_6_out_valid = PE_49_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_17_io_to_pes_6_out_bits = PE_49_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_17_io_to_mem_valid = MemController_17_io_rd_data_valid; // @[pearray.scala 251:29]
  assign PENetwork_17_io_to_mem_bits = MemController_17_io_rd_data_bits; // @[pearray.scala 251:29]
  assign PENetwork_18_io_to_pes_0_out_valid = PE_2_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_18_io_to_pes_0_out_bits = PE_2_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_18_io_to_pes_1_out_valid = PE_10_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_18_io_to_pes_1_out_bits = PE_10_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_18_io_to_pes_2_out_valid = PE_18_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_18_io_to_pes_2_out_bits = PE_18_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_18_io_to_pes_3_out_valid = PE_26_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_18_io_to_pes_3_out_bits = PE_26_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_18_io_to_pes_4_out_valid = PE_34_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_18_io_to_pes_4_out_bits = PE_34_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_18_io_to_pes_5_out_valid = PE_42_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_18_io_to_pes_5_out_bits = PE_42_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_18_io_to_pes_6_out_valid = PE_50_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_18_io_to_pes_6_out_bits = PE_50_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_18_io_to_mem_valid = MemController_18_io_rd_data_valid; // @[pearray.scala 251:29]
  assign PENetwork_18_io_to_mem_bits = MemController_18_io_rd_data_bits; // @[pearray.scala 251:29]
  assign PENetwork_19_io_to_pes_0_out_valid = PE_3_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_19_io_to_pes_0_out_bits = PE_3_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_19_io_to_pes_1_out_valid = PE_11_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_19_io_to_pes_1_out_bits = PE_11_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_19_io_to_pes_2_out_valid = PE_19_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_19_io_to_pes_2_out_bits = PE_19_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_19_io_to_pes_3_out_valid = PE_27_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_19_io_to_pes_3_out_bits = PE_27_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_19_io_to_pes_4_out_valid = PE_35_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_19_io_to_pes_4_out_bits = PE_35_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_19_io_to_pes_5_out_valid = PE_43_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_19_io_to_pes_5_out_bits = PE_43_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_19_io_to_pes_6_out_valid = PE_51_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_19_io_to_pes_6_out_bits = PE_51_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_19_io_to_mem_valid = MemController_19_io_rd_data_valid; // @[pearray.scala 251:29]
  assign PENetwork_19_io_to_mem_bits = MemController_19_io_rd_data_bits; // @[pearray.scala 251:29]
  assign PENetwork_20_io_to_pes_0_out_valid = PE_4_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_20_io_to_pes_0_out_bits = PE_4_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_20_io_to_pes_1_out_valid = PE_12_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_20_io_to_pes_1_out_bits = PE_12_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_20_io_to_pes_2_out_valid = PE_20_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_20_io_to_pes_2_out_bits = PE_20_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_20_io_to_pes_3_out_valid = PE_28_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_20_io_to_pes_3_out_bits = PE_28_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_20_io_to_pes_4_out_valid = PE_36_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_20_io_to_pes_4_out_bits = PE_36_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_20_io_to_pes_5_out_valid = PE_44_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_20_io_to_pes_5_out_bits = PE_44_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_20_io_to_pes_6_out_valid = PE_52_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_20_io_to_pes_6_out_bits = PE_52_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_20_io_to_mem_valid = MemController_20_io_rd_data_valid; // @[pearray.scala 251:29]
  assign PENetwork_20_io_to_mem_bits = MemController_20_io_rd_data_bits; // @[pearray.scala 251:29]
  assign PENetwork_21_io_to_pes_0_out_valid = PE_5_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_21_io_to_pes_0_out_bits = PE_5_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_21_io_to_pes_1_out_valid = PE_13_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_21_io_to_pes_1_out_bits = PE_13_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_21_io_to_pes_2_out_valid = PE_21_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_21_io_to_pes_2_out_bits = PE_21_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_21_io_to_pes_3_out_valid = PE_29_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_21_io_to_pes_3_out_bits = PE_29_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_21_io_to_pes_4_out_valid = PE_37_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_21_io_to_pes_4_out_bits = PE_37_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_21_io_to_pes_5_out_valid = PE_45_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_21_io_to_pes_5_out_bits = PE_45_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_21_io_to_pes_6_out_valid = PE_53_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_21_io_to_pes_6_out_bits = PE_53_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_21_io_to_mem_valid = MemController_21_io_rd_data_valid; // @[pearray.scala 251:29]
  assign PENetwork_21_io_to_mem_bits = MemController_21_io_rd_data_bits; // @[pearray.scala 251:29]
  assign PENetwork_22_io_to_pes_0_out_valid = PE_6_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_22_io_to_pes_0_out_bits = PE_6_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_22_io_to_pes_1_out_valid = PE_14_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_22_io_to_pes_1_out_bits = PE_14_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_22_io_to_pes_2_out_valid = PE_22_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_22_io_to_pes_2_out_bits = PE_22_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_22_io_to_pes_3_out_valid = PE_30_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_22_io_to_pes_3_out_bits = PE_30_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_22_io_to_pes_4_out_valid = PE_38_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_22_io_to_pes_4_out_bits = PE_38_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_22_io_to_pes_5_out_valid = PE_46_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_22_io_to_pes_5_out_bits = PE_46_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_22_io_to_pes_6_out_valid = PE_54_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_22_io_to_pes_6_out_bits = PE_54_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_22_io_to_mem_valid = MemController_22_io_rd_data_valid; // @[pearray.scala 251:29]
  assign PENetwork_22_io_to_mem_bits = MemController_22_io_rd_data_bits; // @[pearray.scala 251:29]
  assign PENetwork_23_io_to_pes_0_out_valid = PE_7_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_23_io_to_pes_0_out_bits = PE_7_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_23_io_to_pes_1_out_valid = PE_15_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_23_io_to_pes_1_out_bits = PE_15_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_23_io_to_pes_2_out_valid = PE_23_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_23_io_to_pes_2_out_bits = PE_23_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_23_io_to_pes_3_out_valid = PE_31_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_23_io_to_pes_3_out_bits = PE_31_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_23_io_to_pes_4_out_valid = PE_39_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_23_io_to_pes_4_out_bits = PE_39_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_23_io_to_pes_5_out_valid = PE_47_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_23_io_to_pes_5_out_bits = PE_47_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_23_io_to_pes_6_out_valid = PE_55_io_data_2_out_valid; // @[pearray.scala 159:36]
  assign PENetwork_23_io_to_pes_6_out_bits = PE_55_io_data_2_out_bits; // @[pearray.scala 159:36]
  assign PENetwork_23_io_to_mem_valid = MemController_23_io_rd_data_valid; // @[pearray.scala 251:29]
  assign PENetwork_23_io_to_mem_bits = MemController_23_io_rd_data_bits; // @[pearray.scala 251:29]
  assign MemController_clock = clock;
  assign MemController_reset = reset;
  assign MemController_io_rd_valid = io_out_valid; // @[pearray.scala 254:28]
  assign MemController_io_wr_valid = PENetwork_io_to_mem_valid; // @[pearray.scala 253:28]
  assign MemController_io_wr_data_valid = PENetwork_io_to_mem_valid; // @[pearray.scala 255:27]
  assign MemController_io_wr_data_bits = PENetwork_io_to_mem_bits; // @[pearray.scala 255:27]
  assign MemController_1_clock = clock;
  assign MemController_1_reset = reset;
  assign MemController_1_io_rd_valid = io_out_valid; // @[pearray.scala 254:28]
  assign MemController_1_io_wr_valid = PENetwork_1_io_to_mem_valid; // @[pearray.scala 253:28]
  assign MemController_1_io_wr_data_valid = PENetwork_1_io_to_mem_valid; // @[pearray.scala 255:27]
  assign MemController_1_io_wr_data_bits = PENetwork_1_io_to_mem_bits; // @[pearray.scala 255:27]
  assign MemController_2_clock = clock;
  assign MemController_2_reset = reset;
  assign MemController_2_io_rd_valid = io_out_valid; // @[pearray.scala 254:28]
  assign MemController_2_io_wr_valid = PENetwork_2_io_to_mem_valid; // @[pearray.scala 253:28]
  assign MemController_2_io_wr_data_valid = PENetwork_2_io_to_mem_valid; // @[pearray.scala 255:27]
  assign MemController_2_io_wr_data_bits = PENetwork_2_io_to_mem_bits; // @[pearray.scala 255:27]
  assign MemController_3_clock = clock;
  assign MemController_3_reset = reset;
  assign MemController_3_io_rd_valid = io_out_valid; // @[pearray.scala 254:28]
  assign MemController_3_io_wr_valid = PENetwork_3_io_to_mem_valid; // @[pearray.scala 253:28]
  assign MemController_3_io_wr_data_valid = PENetwork_3_io_to_mem_valid; // @[pearray.scala 255:27]
  assign MemController_3_io_wr_data_bits = PENetwork_3_io_to_mem_bits; // @[pearray.scala 255:27]
  assign MemController_4_clock = clock;
  assign MemController_4_reset = reset;
  assign MemController_4_io_rd_valid = io_out_valid; // @[pearray.scala 254:28]
  assign MemController_4_io_wr_valid = PENetwork_4_io_to_mem_valid; // @[pearray.scala 253:28]
  assign MemController_4_io_wr_data_valid = PENetwork_4_io_to_mem_valid; // @[pearray.scala 255:27]
  assign MemController_4_io_wr_data_bits = PENetwork_4_io_to_mem_bits; // @[pearray.scala 255:27]
  assign MemController_5_clock = clock;
  assign MemController_5_reset = reset;
  assign MemController_5_io_rd_valid = io_out_valid; // @[pearray.scala 254:28]
  assign MemController_5_io_wr_valid = PENetwork_5_io_to_mem_valid; // @[pearray.scala 253:28]
  assign MemController_5_io_wr_data_valid = PENetwork_5_io_to_mem_valid; // @[pearray.scala 255:27]
  assign MemController_5_io_wr_data_bits = PENetwork_5_io_to_mem_bits; // @[pearray.scala 255:27]
  assign MemController_6_clock = clock;
  assign MemController_6_reset = reset;
  assign MemController_6_io_rd_valid = io_out_valid; // @[pearray.scala 254:28]
  assign MemController_6_io_wr_valid = PENetwork_6_io_to_mem_valid; // @[pearray.scala 253:28]
  assign MemController_6_io_wr_data_valid = PENetwork_6_io_to_mem_valid; // @[pearray.scala 255:27]
  assign MemController_6_io_wr_data_bits = PENetwork_6_io_to_mem_bits; // @[pearray.scala 255:27]
  assign MemController_7_clock = clock;
  assign MemController_7_reset = reset;
  assign MemController_7_io_rd_valid = io_out_valid; // @[pearray.scala 254:28]
  assign MemController_7_io_wr_valid = PENetwork_7_io_to_mem_valid; // @[pearray.scala 253:28]
  assign MemController_7_io_wr_data_valid = PENetwork_7_io_to_mem_valid; // @[pearray.scala 255:27]
  assign MemController_7_io_wr_data_bits = PENetwork_7_io_to_mem_bits; // @[pearray.scala 255:27]
  assign MemController_8_clock = clock;
  assign MemController_8_reset = reset;
  assign MemController_8_io_rd_valid = _T_655_2; // @[pearray.scala 248:30]
  assign MemController_8_io_wr_valid = io_data_1_in_0_valid; // @[pearray.scala 249:28]
  assign MemController_8_io_wr_data_valid = io_data_1_in_0_bits_valid; // @[pearray.scala 250:27]
  assign MemController_8_io_wr_data_bits = io_data_1_in_0_bits_bits; // @[pearray.scala 250:27]
  assign MemController_9_clock = clock;
  assign MemController_9_reset = reset;
  assign MemController_9_io_rd_valid = _T_664_2; // @[pearray.scala 248:30]
  assign MemController_9_io_wr_valid = io_data_1_in_1_valid; // @[pearray.scala 249:28]
  assign MemController_9_io_wr_data_valid = io_data_1_in_1_bits_valid; // @[pearray.scala 250:27]
  assign MemController_9_io_wr_data_bits = io_data_1_in_1_bits_bits; // @[pearray.scala 250:27]
  assign MemController_10_clock = clock;
  assign MemController_10_reset = reset;
  assign MemController_10_io_rd_valid = _T_673_2; // @[pearray.scala 248:30]
  assign MemController_10_io_wr_valid = io_data_1_in_2_valid; // @[pearray.scala 249:28]
  assign MemController_10_io_wr_data_valid = io_data_1_in_2_bits_valid; // @[pearray.scala 250:27]
  assign MemController_10_io_wr_data_bits = io_data_1_in_2_bits_bits; // @[pearray.scala 250:27]
  assign MemController_11_clock = clock;
  assign MemController_11_reset = reset;
  assign MemController_11_io_rd_valid = _T_682_2; // @[pearray.scala 248:30]
  assign MemController_11_io_wr_valid = io_data_1_in_3_valid; // @[pearray.scala 249:28]
  assign MemController_11_io_wr_data_valid = io_data_1_in_3_bits_valid; // @[pearray.scala 250:27]
  assign MemController_11_io_wr_data_bits = io_data_1_in_3_bits_bits; // @[pearray.scala 250:27]
  assign MemController_12_clock = clock;
  assign MemController_12_reset = reset;
  assign MemController_12_io_rd_valid = _T_691_2; // @[pearray.scala 248:30]
  assign MemController_12_io_wr_valid = io_data_1_in_4_valid; // @[pearray.scala 249:28]
  assign MemController_12_io_wr_data_valid = io_data_1_in_4_bits_valid; // @[pearray.scala 250:27]
  assign MemController_12_io_wr_data_bits = io_data_1_in_4_bits_bits; // @[pearray.scala 250:27]
  assign MemController_13_clock = clock;
  assign MemController_13_reset = reset;
  assign MemController_13_io_rd_valid = _T_700_2; // @[pearray.scala 248:30]
  assign MemController_13_io_wr_valid = io_data_1_in_5_valid; // @[pearray.scala 249:28]
  assign MemController_13_io_wr_data_valid = io_data_1_in_5_bits_valid; // @[pearray.scala 250:27]
  assign MemController_13_io_wr_data_bits = io_data_1_in_5_bits_bits; // @[pearray.scala 250:27]
  assign MemController_14_clock = clock;
  assign MemController_14_reset = reset;
  assign MemController_14_io_rd_valid = _T_709_2; // @[pearray.scala 248:30]
  assign MemController_14_io_wr_valid = io_data_1_in_6_valid; // @[pearray.scala 249:28]
  assign MemController_14_io_wr_data_valid = io_data_1_in_6_bits_valid; // @[pearray.scala 250:27]
  assign MemController_14_io_wr_data_bits = io_data_1_in_6_bits_bits; // @[pearray.scala 250:27]
  assign MemController_15_clock = clock;
  assign MemController_15_reset = reset;
  assign MemController_15_io_rd_valid = _T_718_2; // @[pearray.scala 248:30]
  assign MemController_15_io_wr_valid = io_data_1_in_7_valid; // @[pearray.scala 249:28]
  assign MemController_15_io_wr_data_valid = io_data_1_in_7_bits_valid; // @[pearray.scala 250:27]
  assign MemController_15_io_wr_data_bits = io_data_1_in_7_bits_bits; // @[pearray.scala 250:27]
  assign MemController_16_clock = clock;
  assign MemController_16_reset = reset;
  assign MemController_16_io_rd_valid = io_exec_valid; // @[pearray.scala 241:32]
  assign MemController_16_io_wr_valid = io_data_2_in_0_valid; // @[pearray.scala 249:28]
  assign MemController_16_io_wr_data_valid = io_data_2_in_0_bits_valid; // @[pearray.scala 250:27]
  assign MemController_16_io_wr_data_bits = io_data_2_in_0_bits_bits; // @[pearray.scala 250:27]
  assign MemController_17_clock = clock;
  assign MemController_17_reset = reset;
  assign MemController_17_io_rd_valid = _T_720_0; // @[pearray.scala 239:32]
  assign MemController_17_io_wr_valid = io_data_2_in_1_valid; // @[pearray.scala 249:28]
  assign MemController_17_io_wr_data_valid = io_data_2_in_1_bits_valid; // @[pearray.scala 250:27]
  assign MemController_17_io_wr_data_bits = io_data_2_in_1_bits_bits; // @[pearray.scala 250:27]
  assign MemController_18_clock = clock;
  assign MemController_18_reset = reset;
  assign MemController_18_io_rd_valid = _T_720_1; // @[pearray.scala 239:32]
  assign MemController_18_io_wr_valid = io_data_2_in_2_valid; // @[pearray.scala 249:28]
  assign MemController_18_io_wr_data_valid = io_data_2_in_2_bits_valid; // @[pearray.scala 250:27]
  assign MemController_18_io_wr_data_bits = io_data_2_in_2_bits_bits; // @[pearray.scala 250:27]
  assign MemController_19_clock = clock;
  assign MemController_19_reset = reset;
  assign MemController_19_io_rd_valid = _T_720_2; // @[pearray.scala 239:32]
  assign MemController_19_io_wr_valid = io_data_2_in_3_valid; // @[pearray.scala 249:28]
  assign MemController_19_io_wr_data_valid = io_data_2_in_3_bits_valid; // @[pearray.scala 250:27]
  assign MemController_19_io_wr_data_bits = io_data_2_in_3_bits_bits; // @[pearray.scala 250:27]
  assign MemController_20_clock = clock;
  assign MemController_20_reset = reset;
  assign MemController_20_io_rd_valid = _T_720_3; // @[pearray.scala 239:32]
  assign MemController_20_io_wr_valid = io_data_2_in_4_valid; // @[pearray.scala 249:28]
  assign MemController_20_io_wr_data_valid = io_data_2_in_4_bits_valid; // @[pearray.scala 250:27]
  assign MemController_20_io_wr_data_bits = io_data_2_in_4_bits_bits; // @[pearray.scala 250:27]
  assign MemController_21_clock = clock;
  assign MemController_21_reset = reset;
  assign MemController_21_io_rd_valid = _T_720_4; // @[pearray.scala 239:32]
  assign MemController_21_io_wr_valid = io_data_2_in_5_valid; // @[pearray.scala 249:28]
  assign MemController_21_io_wr_data_valid = io_data_2_in_5_bits_valid; // @[pearray.scala 250:27]
  assign MemController_21_io_wr_data_bits = io_data_2_in_5_bits_bits; // @[pearray.scala 250:27]
  assign MemController_22_clock = clock;
  assign MemController_22_reset = reset;
  assign MemController_22_io_rd_valid = _T_720_5; // @[pearray.scala 239:32]
  assign MemController_22_io_wr_valid = io_data_2_in_6_valid; // @[pearray.scala 249:28]
  assign MemController_22_io_wr_data_valid = io_data_2_in_6_bits_valid; // @[pearray.scala 250:27]
  assign MemController_22_io_wr_data_bits = io_data_2_in_6_bits_bits; // @[pearray.scala 250:27]
  assign MemController_23_clock = clock;
  assign MemController_23_reset = reset;
  assign MemController_23_io_rd_valid = _T_720_6; // @[pearray.scala 239:32]
  assign MemController_23_io_wr_valid = io_data_2_in_7_valid; // @[pearray.scala 249:28]
  assign MemController_23_io_wr_data_valid = io_data_2_in_7_bits_valid; // @[pearray.scala 250:27]
  assign MemController_23_io_wr_data_bits = io_data_2_in_7_bits_bits; // @[pearray.scala 250:27]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_12_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_12_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_12_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_12_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_22_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_22_1 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_22_2 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_22_3 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_32_0 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_32_1 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_32_2 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_32_3 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_42_0 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_42_1 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_42_2 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_42_3 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_52_0 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_52_1 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_52_2 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_52_3 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_62_0 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_62_1 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_62_2 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_62_3 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_72_0 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_72_1 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_72_2 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_72_3 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_82_0 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_82_1 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_82_2 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_82_3 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_92_0 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_92_1 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_92_2 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_92_3 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_102_0 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_102_1 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_102_2 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_102_3 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_112_0 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_112_1 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_112_2 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_112_3 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_122_0 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_122_1 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_122_2 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_122_3 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_132_0 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_132_1 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_132_2 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_132_3 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _T_142_0 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _T_142_1 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T_142_2 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T_142_3 = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _T_152_0 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _T_152_1 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T_152_2 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T_152_3 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _T_162_0 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _T_162_1 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T_162_2 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T_162_3 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _T_172_0 = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _T_172_1 = _RAND_65[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _T_172_2 = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _T_172_3 = _RAND_67[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _T_182_0 = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  _T_182_1 = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _T_182_2 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _T_182_3 = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  _T_192_0 = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  _T_192_1 = _RAND_73[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _T_192_2 = _RAND_74[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _T_192_3 = _RAND_75[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  _T_202_0 = _RAND_76[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  _T_202_1 = _RAND_77[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  _T_202_2 = _RAND_78[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  _T_202_3 = _RAND_79[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  _T_212_0 = _RAND_80[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  _T_212_1 = _RAND_81[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _T_212_2 = _RAND_82[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _T_212_3 = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  _T_222_0 = _RAND_84[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  _T_222_1 = _RAND_85[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _T_222_2 = _RAND_86[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  _T_222_3 = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  _T_232_0 = _RAND_88[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  _T_232_1 = _RAND_89[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  _T_232_2 = _RAND_90[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  _T_232_3 = _RAND_91[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  _T_242_0 = _RAND_92[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  _T_242_1 = _RAND_93[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _T_242_2 = _RAND_94[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  _T_242_3 = _RAND_95[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  _T_252_0 = _RAND_96[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  _T_252_1 = _RAND_97[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  _T_252_2 = _RAND_98[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  _T_252_3 = _RAND_99[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  _T_262_0 = _RAND_100[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  _T_262_1 = _RAND_101[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  _T_262_2 = _RAND_102[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  _T_262_3 = _RAND_103[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  _T_272_0 = _RAND_104[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  _T_272_1 = _RAND_105[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  _T_272_2 = _RAND_106[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  _T_272_3 = _RAND_107[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  _T_282_0 = _RAND_108[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  _T_282_1 = _RAND_109[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  _T_282_2 = _RAND_110[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  _T_282_3 = _RAND_111[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  _T_292_0 = _RAND_112[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  _T_292_1 = _RAND_113[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  _T_292_2 = _RAND_114[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  _T_292_3 = _RAND_115[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  _T_302_0 = _RAND_116[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  _T_302_1 = _RAND_117[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  _T_302_2 = _RAND_118[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  _T_302_3 = _RAND_119[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  _T_312_0 = _RAND_120[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  _T_312_1 = _RAND_121[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  _T_312_2 = _RAND_122[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  _T_312_3 = _RAND_123[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  _T_322_0 = _RAND_124[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  _T_322_1 = _RAND_125[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  _T_322_2 = _RAND_126[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  _T_322_3 = _RAND_127[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  _T_332_0 = _RAND_128[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  _T_332_1 = _RAND_129[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  _T_332_2 = _RAND_130[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  _T_332_3 = _RAND_131[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  _T_342_0 = _RAND_132[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  _T_342_1 = _RAND_133[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  _T_342_2 = _RAND_134[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  _T_342_3 = _RAND_135[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  _T_352_0 = _RAND_136[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  _T_352_1 = _RAND_137[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  _T_352_2 = _RAND_138[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  _T_352_3 = _RAND_139[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  _T_362_0 = _RAND_140[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  _T_362_1 = _RAND_141[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  _T_362_2 = _RAND_142[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  _T_362_3 = _RAND_143[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  _T_372_0 = _RAND_144[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  _T_372_1 = _RAND_145[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  _T_372_2 = _RAND_146[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  _T_372_3 = _RAND_147[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  _T_382_0 = _RAND_148[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  _T_382_1 = _RAND_149[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  _T_382_2 = _RAND_150[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  _T_382_3 = _RAND_151[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  _T_392_0 = _RAND_152[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  _T_392_1 = _RAND_153[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  _T_392_2 = _RAND_154[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  _T_392_3 = _RAND_155[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  _T_402_0 = _RAND_156[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  _T_402_1 = _RAND_157[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  _T_402_2 = _RAND_158[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  _T_402_3 = _RAND_159[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  _T_412_0 = _RAND_160[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  _T_412_1 = _RAND_161[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  _T_412_2 = _RAND_162[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  _T_412_3 = _RAND_163[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  _T_422_0 = _RAND_164[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  _T_422_1 = _RAND_165[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  _T_422_2 = _RAND_166[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  _T_422_3 = _RAND_167[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  _T_432_0 = _RAND_168[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  _T_432_1 = _RAND_169[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  _T_432_2 = _RAND_170[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  _T_432_3 = _RAND_171[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  _T_442_0 = _RAND_172[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  _T_442_1 = _RAND_173[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  _T_442_2 = _RAND_174[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  _T_442_3 = _RAND_175[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  _T_452_0 = _RAND_176[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  _T_452_1 = _RAND_177[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  _T_452_2 = _RAND_178[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  _T_452_3 = _RAND_179[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  _T_462_0 = _RAND_180[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  _T_462_1 = _RAND_181[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  _T_462_2 = _RAND_182[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  _T_462_3 = _RAND_183[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  _T_472_0 = _RAND_184[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  _T_472_1 = _RAND_185[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  _T_472_2 = _RAND_186[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  _T_472_3 = _RAND_187[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  _T_482_0 = _RAND_188[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  _T_482_1 = _RAND_189[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  _T_482_2 = _RAND_190[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  _T_482_3 = _RAND_191[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  _T_492_0 = _RAND_192[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  _T_492_1 = _RAND_193[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  _T_492_2 = _RAND_194[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  _T_492_3 = _RAND_195[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  _T_502_0 = _RAND_196[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  _T_502_1 = _RAND_197[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  _T_502_2 = _RAND_198[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  _T_502_3 = _RAND_199[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  _T_512_0 = _RAND_200[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  _T_512_1 = _RAND_201[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  _T_512_2 = _RAND_202[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  _T_512_3 = _RAND_203[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  _T_522_0 = _RAND_204[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  _T_522_1 = _RAND_205[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  _T_522_2 = _RAND_206[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  _T_522_3 = _RAND_207[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  _T_532_0 = _RAND_208[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  _T_532_1 = _RAND_209[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  _T_532_2 = _RAND_210[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  _T_532_3 = _RAND_211[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{`RANDOM}};
  _T_542_0 = _RAND_212[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{`RANDOM}};
  _T_542_1 = _RAND_213[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{`RANDOM}};
  _T_542_2 = _RAND_214[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{`RANDOM}};
  _T_542_3 = _RAND_215[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{`RANDOM}};
  _T_552_0 = _RAND_216[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{`RANDOM}};
  _T_552_1 = _RAND_217[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{`RANDOM}};
  _T_552_2 = _RAND_218[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{`RANDOM}};
  _T_552_3 = _RAND_219[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{`RANDOM}};
  _T_562_0 = _RAND_220[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{`RANDOM}};
  _T_562_1 = _RAND_221[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{`RANDOM}};
  _T_562_2 = _RAND_222[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{`RANDOM}};
  _T_562_3 = _RAND_223[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{`RANDOM}};
  _T_572_0 = _RAND_224[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{`RANDOM}};
  _T_572_1 = _RAND_225[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{`RANDOM}};
  _T_572_2 = _RAND_226[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{`RANDOM}};
  _T_572_3 = _RAND_227[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{`RANDOM}};
  _T_582_0 = _RAND_228[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{`RANDOM}};
  _T_582_1 = _RAND_229[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{`RANDOM}};
  _T_582_2 = _RAND_230[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{`RANDOM}};
  _T_582_3 = _RAND_231[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{`RANDOM}};
  _T_592_0 = _RAND_232[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{`RANDOM}};
  _T_592_1 = _RAND_233[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{`RANDOM}};
  _T_592_2 = _RAND_234[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{`RANDOM}};
  _T_592_3 = _RAND_235[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{`RANDOM}};
  _T_602_0 = _RAND_236[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{`RANDOM}};
  _T_602_1 = _RAND_237[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{`RANDOM}};
  _T_602_2 = _RAND_238[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{`RANDOM}};
  _T_602_3 = _RAND_239[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{`RANDOM}};
  _T_612_0 = _RAND_240[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{`RANDOM}};
  _T_612_1 = _RAND_241[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{`RANDOM}};
  _T_612_2 = _RAND_242[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{`RANDOM}};
  _T_612_3 = _RAND_243[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{`RANDOM}};
  _T_622_0 = _RAND_244[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{`RANDOM}};
  _T_622_1 = _RAND_245[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{`RANDOM}};
  _T_622_2 = _RAND_246[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{`RANDOM}};
  _T_622_3 = _RAND_247[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{`RANDOM}};
  _T_632_0 = _RAND_248[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{`RANDOM}};
  _T_632_1 = _RAND_249[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{`RANDOM}};
  _T_632_2 = _RAND_250[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{`RANDOM}};
  _T_632_3 = _RAND_251[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{`RANDOM}};
  _T_642_0 = _RAND_252[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{`RANDOM}};
  _T_642_1 = _RAND_253[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{`RANDOM}};
  _T_642_2 = _RAND_254[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{`RANDOM}};
  _T_642_3 = _RAND_255[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{`RANDOM}};
  _T_655_0 = _RAND_256[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{`RANDOM}};
  _T_655_1 = _RAND_257[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_258 = {1{`RANDOM}};
  _T_655_2 = _RAND_258[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_259 = {1{`RANDOM}};
  _T_664_0 = _RAND_259[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_260 = {1{`RANDOM}};
  _T_664_1 = _RAND_260[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_261 = {1{`RANDOM}};
  _T_664_2 = _RAND_261[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_262 = {1{`RANDOM}};
  _T_673_0 = _RAND_262[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_263 = {1{`RANDOM}};
  _T_673_1 = _RAND_263[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_264 = {1{`RANDOM}};
  _T_673_2 = _RAND_264[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_265 = {1{`RANDOM}};
  _T_682_0 = _RAND_265[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_266 = {1{`RANDOM}};
  _T_682_1 = _RAND_266[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_267 = {1{`RANDOM}};
  _T_682_2 = _RAND_267[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_268 = {1{`RANDOM}};
  _T_691_0 = _RAND_268[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_269 = {1{`RANDOM}};
  _T_691_1 = _RAND_269[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_270 = {1{`RANDOM}};
  _T_691_2 = _RAND_270[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_271 = {1{`RANDOM}};
  _T_700_0 = _RAND_271[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_272 = {1{`RANDOM}};
  _T_700_1 = _RAND_272[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_273 = {1{`RANDOM}};
  _T_700_2 = _RAND_273[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_274 = {1{`RANDOM}};
  _T_709_0 = _RAND_274[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_275 = {1{`RANDOM}};
  _T_709_1 = _RAND_275[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_276 = {1{`RANDOM}};
  _T_709_2 = _RAND_276[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_277 = {1{`RANDOM}};
  _T_718_0 = _RAND_277[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_278 = {1{`RANDOM}};
  _T_718_1 = _RAND_278[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_279 = {1{`RANDOM}};
  _T_718_2 = _RAND_279[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_280 = {1{`RANDOM}};
  _T_720_0 = _RAND_280[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_281 = {1{`RANDOM}};
  _T_720_1 = _RAND_281[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_282 = {1{`RANDOM}};
  _T_720_2 = _RAND_282[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_283 = {1{`RANDOM}};
  _T_720_3 = _RAND_283[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_284 = {1{`RANDOM}};
  _T_720_4 = _RAND_284[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_285 = {1{`RANDOM}};
  _T_720_5 = _RAND_285[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_286 = {1{`RANDOM}};
  _T_720_6 = _RAND_286[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_12_0 <= 1'h0;
    end else begin
      _T_12_0 <= _T_5;
    end
    if (reset) begin
      _T_12_1 <= 1'h0;
    end else begin
      _T_12_1 <= _T_12_0;
    end
    if (reset) begin
      _T_12_2 <= 1'h0;
    end else begin
      _T_12_2 <= _T_12_1;
    end
    if (reset) begin
      _T_12_3 <= 1'h0;
    end else begin
      _T_12_3 <= _T_12_2;
    end
    if (reset) begin
      _T_22_0 <= 1'h0;
    end else begin
      _T_22_0 <= _T_15;
    end
    if (reset) begin
      _T_22_1 <= 1'h0;
    end else begin
      _T_22_1 <= _T_22_0;
    end
    if (reset) begin
      _T_22_2 <= 1'h0;
    end else begin
      _T_22_2 <= _T_22_1;
    end
    if (reset) begin
      _T_22_3 <= 1'h0;
    end else begin
      _T_22_3 <= _T_22_2;
    end
    if (reset) begin
      _T_32_0 <= 1'h0;
    end else begin
      _T_32_0 <= _T_25;
    end
    if (reset) begin
      _T_32_1 <= 1'h0;
    end else begin
      _T_32_1 <= _T_32_0;
    end
    if (reset) begin
      _T_32_2 <= 1'h0;
    end else begin
      _T_32_2 <= _T_32_1;
    end
    if (reset) begin
      _T_32_3 <= 1'h0;
    end else begin
      _T_32_3 <= _T_32_2;
    end
    if (reset) begin
      _T_42_0 <= 1'h0;
    end else begin
      _T_42_0 <= _T_35;
    end
    if (reset) begin
      _T_42_1 <= 1'h0;
    end else begin
      _T_42_1 <= _T_42_0;
    end
    if (reset) begin
      _T_42_2 <= 1'h0;
    end else begin
      _T_42_2 <= _T_42_1;
    end
    if (reset) begin
      _T_42_3 <= 1'h0;
    end else begin
      _T_42_3 <= _T_42_2;
    end
    if (reset) begin
      _T_52_0 <= 1'h0;
    end else begin
      _T_52_0 <= _T_45;
    end
    if (reset) begin
      _T_52_1 <= 1'h0;
    end else begin
      _T_52_1 <= _T_52_0;
    end
    if (reset) begin
      _T_52_2 <= 1'h0;
    end else begin
      _T_52_2 <= _T_52_1;
    end
    if (reset) begin
      _T_52_3 <= 1'h0;
    end else begin
      _T_52_3 <= _T_52_2;
    end
    if (reset) begin
      _T_62_0 <= 1'h0;
    end else begin
      _T_62_0 <= _T_55;
    end
    if (reset) begin
      _T_62_1 <= 1'h0;
    end else begin
      _T_62_1 <= _T_62_0;
    end
    if (reset) begin
      _T_62_2 <= 1'h0;
    end else begin
      _T_62_2 <= _T_62_1;
    end
    if (reset) begin
      _T_62_3 <= 1'h0;
    end else begin
      _T_62_3 <= _T_62_2;
    end
    if (reset) begin
      _T_72_0 <= 1'h0;
    end else begin
      _T_72_0 <= _T_65;
    end
    if (reset) begin
      _T_72_1 <= 1'h0;
    end else begin
      _T_72_1 <= _T_72_0;
    end
    if (reset) begin
      _T_72_2 <= 1'h0;
    end else begin
      _T_72_2 <= _T_72_1;
    end
    if (reset) begin
      _T_72_3 <= 1'h0;
    end else begin
      _T_72_3 <= _T_72_2;
    end
    if (reset) begin
      _T_82_0 <= 1'h0;
    end else begin
      _T_82_0 <= _T_75;
    end
    if (reset) begin
      _T_82_1 <= 1'h0;
    end else begin
      _T_82_1 <= _T_82_0;
    end
    if (reset) begin
      _T_82_2 <= 1'h0;
    end else begin
      _T_82_2 <= _T_82_1;
    end
    if (reset) begin
      _T_82_3 <= 1'h0;
    end else begin
      _T_82_3 <= _T_82_2;
    end
    if (reset) begin
      _T_92_0 <= 1'h0;
    end else begin
      _T_92_0 <= _T_15;
    end
    if (reset) begin
      _T_92_1 <= 1'h0;
    end else begin
      _T_92_1 <= _T_92_0;
    end
    if (reset) begin
      _T_92_2 <= 1'h0;
    end else begin
      _T_92_2 <= _T_92_1;
    end
    if (reset) begin
      _T_92_3 <= 1'h0;
    end else begin
      _T_92_3 <= _T_92_2;
    end
    if (reset) begin
      _T_102_0 <= 1'h0;
    end else begin
      _T_102_0 <= _T_25;
    end
    if (reset) begin
      _T_102_1 <= 1'h0;
    end else begin
      _T_102_1 <= _T_102_0;
    end
    if (reset) begin
      _T_102_2 <= 1'h0;
    end else begin
      _T_102_2 <= _T_102_1;
    end
    if (reset) begin
      _T_102_3 <= 1'h0;
    end else begin
      _T_102_3 <= _T_102_2;
    end
    if (reset) begin
      _T_112_0 <= 1'h0;
    end else begin
      _T_112_0 <= _T_35;
    end
    if (reset) begin
      _T_112_1 <= 1'h0;
    end else begin
      _T_112_1 <= _T_112_0;
    end
    if (reset) begin
      _T_112_2 <= 1'h0;
    end else begin
      _T_112_2 <= _T_112_1;
    end
    if (reset) begin
      _T_112_3 <= 1'h0;
    end else begin
      _T_112_3 <= _T_112_2;
    end
    if (reset) begin
      _T_122_0 <= 1'h0;
    end else begin
      _T_122_0 <= _T_45;
    end
    if (reset) begin
      _T_122_1 <= 1'h0;
    end else begin
      _T_122_1 <= _T_122_0;
    end
    if (reset) begin
      _T_122_2 <= 1'h0;
    end else begin
      _T_122_2 <= _T_122_1;
    end
    if (reset) begin
      _T_122_3 <= 1'h0;
    end else begin
      _T_122_3 <= _T_122_2;
    end
    if (reset) begin
      _T_132_0 <= 1'h0;
    end else begin
      _T_132_0 <= _T_55;
    end
    if (reset) begin
      _T_132_1 <= 1'h0;
    end else begin
      _T_132_1 <= _T_132_0;
    end
    if (reset) begin
      _T_132_2 <= 1'h0;
    end else begin
      _T_132_2 <= _T_132_1;
    end
    if (reset) begin
      _T_132_3 <= 1'h0;
    end else begin
      _T_132_3 <= _T_132_2;
    end
    if (reset) begin
      _T_142_0 <= 1'h0;
    end else begin
      _T_142_0 <= _T_65;
    end
    if (reset) begin
      _T_142_1 <= 1'h0;
    end else begin
      _T_142_1 <= _T_142_0;
    end
    if (reset) begin
      _T_142_2 <= 1'h0;
    end else begin
      _T_142_2 <= _T_142_1;
    end
    if (reset) begin
      _T_142_3 <= 1'h0;
    end else begin
      _T_142_3 <= _T_142_2;
    end
    if (reset) begin
      _T_152_0 <= 1'h0;
    end else begin
      _T_152_0 <= _T_75;
    end
    if (reset) begin
      _T_152_1 <= 1'h0;
    end else begin
      _T_152_1 <= _T_152_0;
    end
    if (reset) begin
      _T_152_2 <= 1'h0;
    end else begin
      _T_152_2 <= _T_152_1;
    end
    if (reset) begin
      _T_152_3 <= 1'h0;
    end else begin
      _T_152_3 <= _T_152_2;
    end
    if (reset) begin
      _T_162_0 <= 1'h0;
    end else begin
      _T_162_0 <= _T_155;
    end
    if (reset) begin
      _T_162_1 <= 1'h0;
    end else begin
      _T_162_1 <= _T_162_0;
    end
    if (reset) begin
      _T_162_2 <= 1'h0;
    end else begin
      _T_162_2 <= _T_162_1;
    end
    if (reset) begin
      _T_162_3 <= 1'h0;
    end else begin
      _T_162_3 <= _T_162_2;
    end
    if (reset) begin
      _T_172_0 <= 1'h0;
    end else begin
      _T_172_0 <= _T_25;
    end
    if (reset) begin
      _T_172_1 <= 1'h0;
    end else begin
      _T_172_1 <= _T_172_0;
    end
    if (reset) begin
      _T_172_2 <= 1'h0;
    end else begin
      _T_172_2 <= _T_172_1;
    end
    if (reset) begin
      _T_172_3 <= 1'h0;
    end else begin
      _T_172_3 <= _T_172_2;
    end
    if (reset) begin
      _T_182_0 <= 1'h0;
    end else begin
      _T_182_0 <= _T_35;
    end
    if (reset) begin
      _T_182_1 <= 1'h0;
    end else begin
      _T_182_1 <= _T_182_0;
    end
    if (reset) begin
      _T_182_2 <= 1'h0;
    end else begin
      _T_182_2 <= _T_182_1;
    end
    if (reset) begin
      _T_182_3 <= 1'h0;
    end else begin
      _T_182_3 <= _T_182_2;
    end
    if (reset) begin
      _T_192_0 <= 1'h0;
    end else begin
      _T_192_0 <= _T_45;
    end
    if (reset) begin
      _T_192_1 <= 1'h0;
    end else begin
      _T_192_1 <= _T_192_0;
    end
    if (reset) begin
      _T_192_2 <= 1'h0;
    end else begin
      _T_192_2 <= _T_192_1;
    end
    if (reset) begin
      _T_192_3 <= 1'h0;
    end else begin
      _T_192_3 <= _T_192_2;
    end
    if (reset) begin
      _T_202_0 <= 1'h0;
    end else begin
      _T_202_0 <= _T_55;
    end
    if (reset) begin
      _T_202_1 <= 1'h0;
    end else begin
      _T_202_1 <= _T_202_0;
    end
    if (reset) begin
      _T_202_2 <= 1'h0;
    end else begin
      _T_202_2 <= _T_202_1;
    end
    if (reset) begin
      _T_202_3 <= 1'h0;
    end else begin
      _T_202_3 <= _T_202_2;
    end
    if (reset) begin
      _T_212_0 <= 1'h0;
    end else begin
      _T_212_0 <= _T_65;
    end
    if (reset) begin
      _T_212_1 <= 1'h0;
    end else begin
      _T_212_1 <= _T_212_0;
    end
    if (reset) begin
      _T_212_2 <= 1'h0;
    end else begin
      _T_212_2 <= _T_212_1;
    end
    if (reset) begin
      _T_212_3 <= 1'h0;
    end else begin
      _T_212_3 <= _T_212_2;
    end
    if (reset) begin
      _T_222_0 <= 1'h0;
    end else begin
      _T_222_0 <= _T_75;
    end
    if (reset) begin
      _T_222_1 <= 1'h0;
    end else begin
      _T_222_1 <= _T_222_0;
    end
    if (reset) begin
      _T_222_2 <= 1'h0;
    end else begin
      _T_222_2 <= _T_222_1;
    end
    if (reset) begin
      _T_222_3 <= 1'h0;
    end else begin
      _T_222_3 <= _T_222_2;
    end
    if (reset) begin
      _T_232_0 <= 1'h0;
    end else begin
      _T_232_0 <= _T_155;
    end
    if (reset) begin
      _T_232_1 <= 1'h0;
    end else begin
      _T_232_1 <= _T_232_0;
    end
    if (reset) begin
      _T_232_2 <= 1'h0;
    end else begin
      _T_232_2 <= _T_232_1;
    end
    if (reset) begin
      _T_232_3 <= 1'h0;
    end else begin
      _T_232_3 <= _T_232_2;
    end
    if (reset) begin
      _T_242_0 <= 1'h0;
    end else begin
      _T_242_0 <= _T_235;
    end
    if (reset) begin
      _T_242_1 <= 1'h0;
    end else begin
      _T_242_1 <= _T_242_0;
    end
    if (reset) begin
      _T_242_2 <= 1'h0;
    end else begin
      _T_242_2 <= _T_242_1;
    end
    if (reset) begin
      _T_242_3 <= 1'h0;
    end else begin
      _T_242_3 <= _T_242_2;
    end
    if (reset) begin
      _T_252_0 <= 1'h0;
    end else begin
      _T_252_0 <= _T_35;
    end
    if (reset) begin
      _T_252_1 <= 1'h0;
    end else begin
      _T_252_1 <= _T_252_0;
    end
    if (reset) begin
      _T_252_2 <= 1'h0;
    end else begin
      _T_252_2 <= _T_252_1;
    end
    if (reset) begin
      _T_252_3 <= 1'h0;
    end else begin
      _T_252_3 <= _T_252_2;
    end
    if (reset) begin
      _T_262_0 <= 1'h0;
    end else begin
      _T_262_0 <= _T_45;
    end
    if (reset) begin
      _T_262_1 <= 1'h0;
    end else begin
      _T_262_1 <= _T_262_0;
    end
    if (reset) begin
      _T_262_2 <= 1'h0;
    end else begin
      _T_262_2 <= _T_262_1;
    end
    if (reset) begin
      _T_262_3 <= 1'h0;
    end else begin
      _T_262_3 <= _T_262_2;
    end
    if (reset) begin
      _T_272_0 <= 1'h0;
    end else begin
      _T_272_0 <= _T_55;
    end
    if (reset) begin
      _T_272_1 <= 1'h0;
    end else begin
      _T_272_1 <= _T_272_0;
    end
    if (reset) begin
      _T_272_2 <= 1'h0;
    end else begin
      _T_272_2 <= _T_272_1;
    end
    if (reset) begin
      _T_272_3 <= 1'h0;
    end else begin
      _T_272_3 <= _T_272_2;
    end
    if (reset) begin
      _T_282_0 <= 1'h0;
    end else begin
      _T_282_0 <= _T_65;
    end
    if (reset) begin
      _T_282_1 <= 1'h0;
    end else begin
      _T_282_1 <= _T_282_0;
    end
    if (reset) begin
      _T_282_2 <= 1'h0;
    end else begin
      _T_282_2 <= _T_282_1;
    end
    if (reset) begin
      _T_282_3 <= 1'h0;
    end else begin
      _T_282_3 <= _T_282_2;
    end
    if (reset) begin
      _T_292_0 <= 1'h0;
    end else begin
      _T_292_0 <= _T_75;
    end
    if (reset) begin
      _T_292_1 <= 1'h0;
    end else begin
      _T_292_1 <= _T_292_0;
    end
    if (reset) begin
      _T_292_2 <= 1'h0;
    end else begin
      _T_292_2 <= _T_292_1;
    end
    if (reset) begin
      _T_292_3 <= 1'h0;
    end else begin
      _T_292_3 <= _T_292_2;
    end
    if (reset) begin
      _T_302_0 <= 1'h0;
    end else begin
      _T_302_0 <= _T_155;
    end
    if (reset) begin
      _T_302_1 <= 1'h0;
    end else begin
      _T_302_1 <= _T_302_0;
    end
    if (reset) begin
      _T_302_2 <= 1'h0;
    end else begin
      _T_302_2 <= _T_302_1;
    end
    if (reset) begin
      _T_302_3 <= 1'h0;
    end else begin
      _T_302_3 <= _T_302_2;
    end
    if (reset) begin
      _T_312_0 <= 1'h0;
    end else begin
      _T_312_0 <= _T_235;
    end
    if (reset) begin
      _T_312_1 <= 1'h0;
    end else begin
      _T_312_1 <= _T_312_0;
    end
    if (reset) begin
      _T_312_2 <= 1'h0;
    end else begin
      _T_312_2 <= _T_312_1;
    end
    if (reset) begin
      _T_312_3 <= 1'h0;
    end else begin
      _T_312_3 <= _T_312_2;
    end
    if (reset) begin
      _T_322_0 <= 1'h0;
    end else begin
      _T_322_0 <= _T_315;
    end
    if (reset) begin
      _T_322_1 <= 1'h0;
    end else begin
      _T_322_1 <= _T_322_0;
    end
    if (reset) begin
      _T_322_2 <= 1'h0;
    end else begin
      _T_322_2 <= _T_322_1;
    end
    if (reset) begin
      _T_322_3 <= 1'h0;
    end else begin
      _T_322_3 <= _T_322_2;
    end
    if (reset) begin
      _T_332_0 <= 1'h0;
    end else begin
      _T_332_0 <= _T_45;
    end
    if (reset) begin
      _T_332_1 <= 1'h0;
    end else begin
      _T_332_1 <= _T_332_0;
    end
    if (reset) begin
      _T_332_2 <= 1'h0;
    end else begin
      _T_332_2 <= _T_332_1;
    end
    if (reset) begin
      _T_332_3 <= 1'h0;
    end else begin
      _T_332_3 <= _T_332_2;
    end
    if (reset) begin
      _T_342_0 <= 1'h0;
    end else begin
      _T_342_0 <= _T_55;
    end
    if (reset) begin
      _T_342_1 <= 1'h0;
    end else begin
      _T_342_1 <= _T_342_0;
    end
    if (reset) begin
      _T_342_2 <= 1'h0;
    end else begin
      _T_342_2 <= _T_342_1;
    end
    if (reset) begin
      _T_342_3 <= 1'h0;
    end else begin
      _T_342_3 <= _T_342_2;
    end
    if (reset) begin
      _T_352_0 <= 1'h0;
    end else begin
      _T_352_0 <= _T_65;
    end
    if (reset) begin
      _T_352_1 <= 1'h0;
    end else begin
      _T_352_1 <= _T_352_0;
    end
    if (reset) begin
      _T_352_2 <= 1'h0;
    end else begin
      _T_352_2 <= _T_352_1;
    end
    if (reset) begin
      _T_352_3 <= 1'h0;
    end else begin
      _T_352_3 <= _T_352_2;
    end
    if (reset) begin
      _T_362_0 <= 1'h0;
    end else begin
      _T_362_0 <= _T_75;
    end
    if (reset) begin
      _T_362_1 <= 1'h0;
    end else begin
      _T_362_1 <= _T_362_0;
    end
    if (reset) begin
      _T_362_2 <= 1'h0;
    end else begin
      _T_362_2 <= _T_362_1;
    end
    if (reset) begin
      _T_362_3 <= 1'h0;
    end else begin
      _T_362_3 <= _T_362_2;
    end
    if (reset) begin
      _T_372_0 <= 1'h0;
    end else begin
      _T_372_0 <= _T_155;
    end
    if (reset) begin
      _T_372_1 <= 1'h0;
    end else begin
      _T_372_1 <= _T_372_0;
    end
    if (reset) begin
      _T_372_2 <= 1'h0;
    end else begin
      _T_372_2 <= _T_372_1;
    end
    if (reset) begin
      _T_372_3 <= 1'h0;
    end else begin
      _T_372_3 <= _T_372_2;
    end
    if (reset) begin
      _T_382_0 <= 1'h0;
    end else begin
      _T_382_0 <= _T_235;
    end
    if (reset) begin
      _T_382_1 <= 1'h0;
    end else begin
      _T_382_1 <= _T_382_0;
    end
    if (reset) begin
      _T_382_2 <= 1'h0;
    end else begin
      _T_382_2 <= _T_382_1;
    end
    if (reset) begin
      _T_382_3 <= 1'h0;
    end else begin
      _T_382_3 <= _T_382_2;
    end
    if (reset) begin
      _T_392_0 <= 1'h0;
    end else begin
      _T_392_0 <= _T_315;
    end
    if (reset) begin
      _T_392_1 <= 1'h0;
    end else begin
      _T_392_1 <= _T_392_0;
    end
    if (reset) begin
      _T_392_2 <= 1'h0;
    end else begin
      _T_392_2 <= _T_392_1;
    end
    if (reset) begin
      _T_392_3 <= 1'h0;
    end else begin
      _T_392_3 <= _T_392_2;
    end
    if (reset) begin
      _T_402_0 <= 1'h0;
    end else begin
      _T_402_0 <= _T_395;
    end
    if (reset) begin
      _T_402_1 <= 1'h0;
    end else begin
      _T_402_1 <= _T_402_0;
    end
    if (reset) begin
      _T_402_2 <= 1'h0;
    end else begin
      _T_402_2 <= _T_402_1;
    end
    if (reset) begin
      _T_402_3 <= 1'h0;
    end else begin
      _T_402_3 <= _T_402_2;
    end
    if (reset) begin
      _T_412_0 <= 1'h0;
    end else begin
      _T_412_0 <= _T_55;
    end
    if (reset) begin
      _T_412_1 <= 1'h0;
    end else begin
      _T_412_1 <= _T_412_0;
    end
    if (reset) begin
      _T_412_2 <= 1'h0;
    end else begin
      _T_412_2 <= _T_412_1;
    end
    if (reset) begin
      _T_412_3 <= 1'h0;
    end else begin
      _T_412_3 <= _T_412_2;
    end
    if (reset) begin
      _T_422_0 <= 1'h0;
    end else begin
      _T_422_0 <= _T_65;
    end
    if (reset) begin
      _T_422_1 <= 1'h0;
    end else begin
      _T_422_1 <= _T_422_0;
    end
    if (reset) begin
      _T_422_2 <= 1'h0;
    end else begin
      _T_422_2 <= _T_422_1;
    end
    if (reset) begin
      _T_422_3 <= 1'h0;
    end else begin
      _T_422_3 <= _T_422_2;
    end
    if (reset) begin
      _T_432_0 <= 1'h0;
    end else begin
      _T_432_0 <= _T_75;
    end
    if (reset) begin
      _T_432_1 <= 1'h0;
    end else begin
      _T_432_1 <= _T_432_0;
    end
    if (reset) begin
      _T_432_2 <= 1'h0;
    end else begin
      _T_432_2 <= _T_432_1;
    end
    if (reset) begin
      _T_432_3 <= 1'h0;
    end else begin
      _T_432_3 <= _T_432_2;
    end
    if (reset) begin
      _T_442_0 <= 1'h0;
    end else begin
      _T_442_0 <= _T_155;
    end
    if (reset) begin
      _T_442_1 <= 1'h0;
    end else begin
      _T_442_1 <= _T_442_0;
    end
    if (reset) begin
      _T_442_2 <= 1'h0;
    end else begin
      _T_442_2 <= _T_442_1;
    end
    if (reset) begin
      _T_442_3 <= 1'h0;
    end else begin
      _T_442_3 <= _T_442_2;
    end
    if (reset) begin
      _T_452_0 <= 1'h0;
    end else begin
      _T_452_0 <= _T_235;
    end
    if (reset) begin
      _T_452_1 <= 1'h0;
    end else begin
      _T_452_1 <= _T_452_0;
    end
    if (reset) begin
      _T_452_2 <= 1'h0;
    end else begin
      _T_452_2 <= _T_452_1;
    end
    if (reset) begin
      _T_452_3 <= 1'h0;
    end else begin
      _T_452_3 <= _T_452_2;
    end
    if (reset) begin
      _T_462_0 <= 1'h0;
    end else begin
      _T_462_0 <= _T_315;
    end
    if (reset) begin
      _T_462_1 <= 1'h0;
    end else begin
      _T_462_1 <= _T_462_0;
    end
    if (reset) begin
      _T_462_2 <= 1'h0;
    end else begin
      _T_462_2 <= _T_462_1;
    end
    if (reset) begin
      _T_462_3 <= 1'h0;
    end else begin
      _T_462_3 <= _T_462_2;
    end
    if (reset) begin
      _T_472_0 <= 1'h0;
    end else begin
      _T_472_0 <= _T_395;
    end
    if (reset) begin
      _T_472_1 <= 1'h0;
    end else begin
      _T_472_1 <= _T_472_0;
    end
    if (reset) begin
      _T_472_2 <= 1'h0;
    end else begin
      _T_472_2 <= _T_472_1;
    end
    if (reset) begin
      _T_472_3 <= 1'h0;
    end else begin
      _T_472_3 <= _T_472_2;
    end
    if (reset) begin
      _T_482_0 <= 1'h0;
    end else begin
      _T_482_0 <= _T_475;
    end
    if (reset) begin
      _T_482_1 <= 1'h0;
    end else begin
      _T_482_1 <= _T_482_0;
    end
    if (reset) begin
      _T_482_2 <= 1'h0;
    end else begin
      _T_482_2 <= _T_482_1;
    end
    if (reset) begin
      _T_482_3 <= 1'h0;
    end else begin
      _T_482_3 <= _T_482_2;
    end
    if (reset) begin
      _T_492_0 <= 1'h0;
    end else begin
      _T_492_0 <= _T_65;
    end
    if (reset) begin
      _T_492_1 <= 1'h0;
    end else begin
      _T_492_1 <= _T_492_0;
    end
    if (reset) begin
      _T_492_2 <= 1'h0;
    end else begin
      _T_492_2 <= _T_492_1;
    end
    if (reset) begin
      _T_492_3 <= 1'h0;
    end else begin
      _T_492_3 <= _T_492_2;
    end
    if (reset) begin
      _T_502_0 <= 1'h0;
    end else begin
      _T_502_0 <= _T_75;
    end
    if (reset) begin
      _T_502_1 <= 1'h0;
    end else begin
      _T_502_1 <= _T_502_0;
    end
    if (reset) begin
      _T_502_2 <= 1'h0;
    end else begin
      _T_502_2 <= _T_502_1;
    end
    if (reset) begin
      _T_502_3 <= 1'h0;
    end else begin
      _T_502_3 <= _T_502_2;
    end
    if (reset) begin
      _T_512_0 <= 1'h0;
    end else begin
      _T_512_0 <= _T_155;
    end
    if (reset) begin
      _T_512_1 <= 1'h0;
    end else begin
      _T_512_1 <= _T_512_0;
    end
    if (reset) begin
      _T_512_2 <= 1'h0;
    end else begin
      _T_512_2 <= _T_512_1;
    end
    if (reset) begin
      _T_512_3 <= 1'h0;
    end else begin
      _T_512_3 <= _T_512_2;
    end
    if (reset) begin
      _T_522_0 <= 1'h0;
    end else begin
      _T_522_0 <= _T_235;
    end
    if (reset) begin
      _T_522_1 <= 1'h0;
    end else begin
      _T_522_1 <= _T_522_0;
    end
    if (reset) begin
      _T_522_2 <= 1'h0;
    end else begin
      _T_522_2 <= _T_522_1;
    end
    if (reset) begin
      _T_522_3 <= 1'h0;
    end else begin
      _T_522_3 <= _T_522_2;
    end
    if (reset) begin
      _T_532_0 <= 1'h0;
    end else begin
      _T_532_0 <= _T_315;
    end
    if (reset) begin
      _T_532_1 <= 1'h0;
    end else begin
      _T_532_1 <= _T_532_0;
    end
    if (reset) begin
      _T_532_2 <= 1'h0;
    end else begin
      _T_532_2 <= _T_532_1;
    end
    if (reset) begin
      _T_532_3 <= 1'h0;
    end else begin
      _T_532_3 <= _T_532_2;
    end
    if (reset) begin
      _T_542_0 <= 1'h0;
    end else begin
      _T_542_0 <= _T_395;
    end
    if (reset) begin
      _T_542_1 <= 1'h0;
    end else begin
      _T_542_1 <= _T_542_0;
    end
    if (reset) begin
      _T_542_2 <= 1'h0;
    end else begin
      _T_542_2 <= _T_542_1;
    end
    if (reset) begin
      _T_542_3 <= 1'h0;
    end else begin
      _T_542_3 <= _T_542_2;
    end
    if (reset) begin
      _T_552_0 <= 1'h0;
    end else begin
      _T_552_0 <= _T_475;
    end
    if (reset) begin
      _T_552_1 <= 1'h0;
    end else begin
      _T_552_1 <= _T_552_0;
    end
    if (reset) begin
      _T_552_2 <= 1'h0;
    end else begin
      _T_552_2 <= _T_552_1;
    end
    if (reset) begin
      _T_552_3 <= 1'h0;
    end else begin
      _T_552_3 <= _T_552_2;
    end
    if (reset) begin
      _T_562_0 <= 1'h0;
    end else begin
      _T_562_0 <= _T_555;
    end
    if (reset) begin
      _T_562_1 <= 1'h0;
    end else begin
      _T_562_1 <= _T_562_0;
    end
    if (reset) begin
      _T_562_2 <= 1'h0;
    end else begin
      _T_562_2 <= _T_562_1;
    end
    if (reset) begin
      _T_562_3 <= 1'h0;
    end else begin
      _T_562_3 <= _T_562_2;
    end
    if (reset) begin
      _T_572_0 <= 1'h0;
    end else begin
      _T_572_0 <= _T_75;
    end
    if (reset) begin
      _T_572_1 <= 1'h0;
    end else begin
      _T_572_1 <= _T_572_0;
    end
    if (reset) begin
      _T_572_2 <= 1'h0;
    end else begin
      _T_572_2 <= _T_572_1;
    end
    if (reset) begin
      _T_572_3 <= 1'h0;
    end else begin
      _T_572_3 <= _T_572_2;
    end
    if (reset) begin
      _T_582_0 <= 1'h0;
    end else begin
      _T_582_0 <= _T_155;
    end
    if (reset) begin
      _T_582_1 <= 1'h0;
    end else begin
      _T_582_1 <= _T_582_0;
    end
    if (reset) begin
      _T_582_2 <= 1'h0;
    end else begin
      _T_582_2 <= _T_582_1;
    end
    if (reset) begin
      _T_582_3 <= 1'h0;
    end else begin
      _T_582_3 <= _T_582_2;
    end
    if (reset) begin
      _T_592_0 <= 1'h0;
    end else begin
      _T_592_0 <= _T_235;
    end
    if (reset) begin
      _T_592_1 <= 1'h0;
    end else begin
      _T_592_1 <= _T_592_0;
    end
    if (reset) begin
      _T_592_2 <= 1'h0;
    end else begin
      _T_592_2 <= _T_592_1;
    end
    if (reset) begin
      _T_592_3 <= 1'h0;
    end else begin
      _T_592_3 <= _T_592_2;
    end
    if (reset) begin
      _T_602_0 <= 1'h0;
    end else begin
      _T_602_0 <= _T_315;
    end
    if (reset) begin
      _T_602_1 <= 1'h0;
    end else begin
      _T_602_1 <= _T_602_0;
    end
    if (reset) begin
      _T_602_2 <= 1'h0;
    end else begin
      _T_602_2 <= _T_602_1;
    end
    if (reset) begin
      _T_602_3 <= 1'h0;
    end else begin
      _T_602_3 <= _T_602_2;
    end
    if (reset) begin
      _T_612_0 <= 1'h0;
    end else begin
      _T_612_0 <= _T_395;
    end
    if (reset) begin
      _T_612_1 <= 1'h0;
    end else begin
      _T_612_1 <= _T_612_0;
    end
    if (reset) begin
      _T_612_2 <= 1'h0;
    end else begin
      _T_612_2 <= _T_612_1;
    end
    if (reset) begin
      _T_612_3 <= 1'h0;
    end else begin
      _T_612_3 <= _T_612_2;
    end
    if (reset) begin
      _T_622_0 <= 1'h0;
    end else begin
      _T_622_0 <= _T_475;
    end
    if (reset) begin
      _T_622_1 <= 1'h0;
    end else begin
      _T_622_1 <= _T_622_0;
    end
    if (reset) begin
      _T_622_2 <= 1'h0;
    end else begin
      _T_622_2 <= _T_622_1;
    end
    if (reset) begin
      _T_622_3 <= 1'h0;
    end else begin
      _T_622_3 <= _T_622_2;
    end
    if (reset) begin
      _T_632_0 <= 1'h0;
    end else begin
      _T_632_0 <= _T_555;
    end
    if (reset) begin
      _T_632_1 <= 1'h0;
    end else begin
      _T_632_1 <= _T_632_0;
    end
    if (reset) begin
      _T_632_2 <= 1'h0;
    end else begin
      _T_632_2 <= _T_632_1;
    end
    if (reset) begin
      _T_632_3 <= 1'h0;
    end else begin
      _T_632_3 <= _T_632_2;
    end
    if (reset) begin
      _T_642_0 <= 1'h0;
    end else begin
      _T_642_0 <= _T_635;
    end
    if (reset) begin
      _T_642_1 <= 1'h0;
    end else begin
      _T_642_1 <= _T_642_0;
    end
    if (reset) begin
      _T_642_2 <= 1'h0;
    end else begin
      _T_642_2 <= _T_642_1;
    end
    if (reset) begin
      _T_642_3 <= 1'h0;
    end else begin
      _T_642_3 <= _T_642_2;
    end
    if (reset) begin
      _T_655_0 <= 1'h0;
    end else begin
      _T_655_0 <= _T_650;
    end
    if (reset) begin
      _T_655_1 <= 1'h0;
    end else begin
      _T_655_1 <= _T_655_0;
    end
    if (reset) begin
      _T_655_2 <= 1'h0;
    end else begin
      _T_655_2 <= _T_655_1;
    end
    if (reset) begin
      _T_664_0 <= 1'h0;
    end else begin
      _T_664_0 <= _T_659;
    end
    if (reset) begin
      _T_664_1 <= 1'h0;
    end else begin
      _T_664_1 <= _T_664_0;
    end
    if (reset) begin
      _T_664_2 <= 1'h0;
    end else begin
      _T_664_2 <= _T_664_1;
    end
    if (reset) begin
      _T_673_0 <= 1'h0;
    end else begin
      _T_673_0 <= _T_668;
    end
    if (reset) begin
      _T_673_1 <= 1'h0;
    end else begin
      _T_673_1 <= _T_673_0;
    end
    if (reset) begin
      _T_673_2 <= 1'h0;
    end else begin
      _T_673_2 <= _T_673_1;
    end
    if (reset) begin
      _T_682_0 <= 1'h0;
    end else begin
      _T_682_0 <= _T_677;
    end
    if (reset) begin
      _T_682_1 <= 1'h0;
    end else begin
      _T_682_1 <= _T_682_0;
    end
    if (reset) begin
      _T_682_2 <= 1'h0;
    end else begin
      _T_682_2 <= _T_682_1;
    end
    if (reset) begin
      _T_691_0 <= 1'h0;
    end else begin
      _T_691_0 <= _T_686;
    end
    if (reset) begin
      _T_691_1 <= 1'h0;
    end else begin
      _T_691_1 <= _T_691_0;
    end
    if (reset) begin
      _T_691_2 <= 1'h0;
    end else begin
      _T_691_2 <= _T_691_1;
    end
    if (reset) begin
      _T_700_0 <= 1'h0;
    end else begin
      _T_700_0 <= _T_695;
    end
    if (reset) begin
      _T_700_1 <= 1'h0;
    end else begin
      _T_700_1 <= _T_700_0;
    end
    if (reset) begin
      _T_700_2 <= 1'h0;
    end else begin
      _T_700_2 <= _T_700_1;
    end
    if (reset) begin
      _T_709_0 <= 1'h0;
    end else begin
      _T_709_0 <= _T_704;
    end
    if (reset) begin
      _T_709_1 <= 1'h0;
    end else begin
      _T_709_1 <= _T_709_0;
    end
    if (reset) begin
      _T_709_2 <= 1'h0;
    end else begin
      _T_709_2 <= _T_709_1;
    end
    if (reset) begin
      _T_718_0 <= 1'h0;
    end else begin
      _T_718_0 <= _T_713;
    end
    if (reset) begin
      _T_718_1 <= 1'h0;
    end else begin
      _T_718_1 <= _T_718_0;
    end
    if (reset) begin
      _T_718_2 <= 1'h0;
    end else begin
      _T_718_2 <= _T_718_1;
    end
    if (reset) begin
      _T_720_0 <= 1'h0;
    end else begin
      _T_720_0 <= io_exec_valid;
    end
    if (reset) begin
      _T_720_1 <= 1'h0;
    end else begin
      _T_720_1 <= _T_720_0;
    end
    if (reset) begin
      _T_720_2 <= 1'h0;
    end else begin
      _T_720_2 <= _T_720_1;
    end
    if (reset) begin
      _T_720_3 <= 1'h0;
    end else begin
      _T_720_3 <= _T_720_2;
    end
    if (reset) begin
      _T_720_4 <= 1'h0;
    end else begin
      _T_720_4 <= _T_720_3;
    end
    if (reset) begin
      _T_720_5 <= 1'h0;
    end else begin
      _T_720_5 <= _T_720_4;
    end
    if (reset) begin
      _T_720_6 <= 1'h0;
    end else begin
      _T_720_6 <= _T_720_5;
    end
  end
endmodule
